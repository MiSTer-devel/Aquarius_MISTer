library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity main_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of main_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"E1",X"1F",X"82",X"06",X"22",X"0B",X"00",X"7E",X"E3",X"BE",X"23",X"E3",X"C2",X"C4",X"03",
		X"23",X"7E",X"FE",X"3A",X"D0",X"C3",X"70",X"06",X"C3",X"8A",X"19",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"92",X"C0",X"7D",X"93",X"C9",X"00",X"00",X"3A",X"E7",X"38",X"B7",X"C2",X"EB",X"14",X"C9",
		X"DD",X"2A",X"06",X"38",X"DD",X"E9",X"00",X"00",X"C3",X"03",X"38",X"D9",X"E1",X"23",X"E5",X"D9",
		X"C9",X"31",X"A0",X"38",X"3E",X"0B",X"CD",X"94",X"1D",X"2A",X"01",X"38",X"36",X"20",X"3E",X"07",
		X"CD",X"94",X"1D",X"AF",X"D3",X"FF",X"21",X"FF",X"2F",X"22",X"5D",X"38",X"11",X"11",X"E0",X"21",
		X"81",X"00",X"1B",X"1B",X"23",X"1A",X"0F",X"0F",X"83",X"BE",X"28",X"F6",X"7E",X"B7",X"20",X"19",
		X"EB",X"06",X"0C",X"86",X"23",X"80",X"05",X"20",X"FA",X"AE",X"D3",X"FF",X"32",X"09",X"38",X"C3",
		X"10",X"E0",X"2B",X"37",X"24",X"24",X"33",X"2C",X"00",X"11",X"A1",X"31",X"21",X"B0",X"00",X"01",
		X"05",X"00",X"ED",X"B0",X"11",X"10",X"32",X"21",X"B5",X"00",X"01",X"19",X"00",X"ED",X"B0",X"06",
		X"03",X"CD",X"CF",X"00",X"06",X"02",X"CD",X"CF",X"00",X"06",X"06",X"CD",X"CF",X"00",X"18",X"EF",
		X"42",X"41",X"53",X"49",X"43",X"50",X"72",X"65",X"73",X"73",X"20",X"52",X"45",X"54",X"55",X"52",
		X"4E",X"20",X"6B",X"65",X"79",X"20",X"74",X"6F",X"20",X"73",X"74",X"61",X"72",X"74",X"00",X"21",
		X"00",X"34",X"70",X"23",X"7C",X"FE",X"38",X"20",X"F9",X"21",X"00",X"40",X"CD",X"80",X"1E",X"FE",
		X"0D",X"28",X"1A",X"FE",X"03",X"28",X"06",X"2B",X"7C",X"B5",X"20",X"F0",X"C9",X"3E",X"0B",X"CD",
		X"72",X"1D",X"3A",X"09",X"38",X"D3",X"FF",X"CD",X"E5",X"0B",X"CD",X"40",X"1A",X"21",X"87",X"01",
		X"01",X"51",X"00",X"11",X"03",X"38",X"ED",X"B0",X"AF",X"32",X"A9",X"38",X"32",X"00",X"39",X"21",
		X"64",X"39",X"23",X"4E",X"7C",X"B5",X"28",X"0B",X"A9",X"77",X"46",X"2F",X"77",X"7E",X"2F",X"71",
		X"B8",X"28",X"EF",X"2B",X"11",X"2C",X"3A",X"E7",X"DA",X"B7",X"0B",X"11",X"CE",X"FF",X"22",X"AD",
		X"38",X"19",X"22",X"4B",X"38",X"CD",X"BE",X"0B",X"CD",X"F2",X"1F",X"31",X"65",X"38",X"CD",X"E5",
		X"0B",X"21",X"05",X"20",X"11",X"82",X"00",X"1A",X"B7",X"CA",X"E8",X"1F",X"BE",X"20",X"04",X"2B",
		X"13",X"18",X"F4",X"ED",X"5F",X"17",X"81",X"D3",X"FF",X"32",X"09",X"38",X"C3",X"02",X"04",X"0B",
		X"43",X"6F",X"70",X"79",X"72",X"69",X"67",X"68",X"74",X"20",X"05",X"20",X"31",X"39",X"38",X"32",
		X"20",X"62",X"79",X"20",X"4D",X"69",X"63",X"72",X"6F",X"73",X"6F",X"66",X"74",X"20",X"49",X"6E",
		X"63",X"2E",X"20",X"53",X"32",X"0A",X"00",X"C3",X"97",X"06",X"3B",X"00",X"00",X"A3",X"00",X"00",
		X"00",X"20",X"00",X"00",X"D6",X"00",X"6F",X"7C",X"DE",X"00",X"67",X"78",X"DE",X"00",X"47",X"3E",
		X"00",X"C9",X"00",X"00",X"00",X"35",X"4A",X"CA",X"99",X"39",X"1C",X"76",X"98",X"22",X"95",X"B3",
		X"98",X"0A",X"DD",X"47",X"98",X"53",X"D1",X"99",X"99",X"0A",X"1A",X"9F",X"98",X"65",X"BC",X"CD",
		X"98",X"D6",X"77",X"3E",X"98",X"52",X"C7",X"4F",X"80",X"00",X"00",X"00",X"28",X"0E",X"00",X"64",
		X"39",X"FE",X"FF",X"01",X"39",X"21",X"0C",X"BC",X"05",X"13",X"0D",X"1C",X"07",X"93",X"08",X"CC",
		X"10",X"BE",X"08",X"31",X"07",X"DC",X"06",X"BE",X"06",X"9C",X"07",X"05",X"0C",X"CB",X"06",X"F8",
		X"06",X"1E",X"07",X"1F",X"0C",X"80",X"07",X"B5",X"07",X"15",X"1B",X"3B",X"0B",X"6D",X"0B",X"BC",
		X"07",X"4B",X"0C",X"6C",X"05",X"67",X"05",X"CD",X"0C",X"2C",X"1C",X"08",X"1C",X"4F",X"1A",X"4C",
		X"1A",X"D6",X"1A",X"BD",X"0B",X"F5",X"14",X"B1",X"15",X"09",X"15",X"03",X"38",X"A8",X"10",X"2E",
		X"0B",X"33",X"0B",X"75",X"17",X"66",X"18",X"85",X"13",X"CD",X"17",X"D7",X"18",X"DD",X"18",X"70",
		X"19",X"85",X"19",X"63",X"0B",X"F3",X"0F",X"29",X"0E",X"84",X"10",X"02",X"10",X"13",X"10",X"21",
		X"10",X"50",X"10",X"59",X"10",X"C5",X"4E",X"44",X"C6",X"4F",X"52",X"CE",X"45",X"58",X"54",X"C4",
		X"41",X"54",X"41",X"C9",X"4E",X"50",X"55",X"54",X"C4",X"49",X"4D",X"D2",X"45",X"41",X"44",X"CC",
		X"45",X"54",X"C7",X"4F",X"54",X"4F",X"D2",X"55",X"4E",X"C9",X"46",X"D2",X"45",X"53",X"54",X"4F",
		X"52",X"45",X"C7",X"4F",X"53",X"55",X"42",X"D2",X"45",X"54",X"55",X"52",X"4E",X"D2",X"45",X"4D",
		X"D3",X"54",X"4F",X"50",X"CF",X"4E",X"CC",X"50",X"52",X"49",X"4E",X"54",X"C3",X"4F",X"50",X"59",
		X"C4",X"45",X"46",X"D0",X"4F",X"4B",X"45",X"D0",X"52",X"49",X"4E",X"54",X"C3",X"4F",X"4E",X"54",
		X"CC",X"49",X"53",X"54",X"CC",X"4C",X"49",X"53",X"54",X"C3",X"4C",X"45",X"41",X"52",X"C3",X"4C",
		X"4F",X"41",X"44",X"C3",X"53",X"41",X"56",X"45",X"D0",X"53",X"45",X"54",X"D0",X"52",X"45",X"53",
		X"45",X"54",X"D3",X"4F",X"55",X"4E",X"44",X"CE",X"45",X"57",X"D4",X"41",X"42",X"28",X"D4",X"4F",
		X"C6",X"4E",X"D3",X"50",X"43",X"28",X"C9",X"4E",X"4B",X"45",X"59",X"24",X"D4",X"48",X"45",X"4E",
		X"CE",X"4F",X"54",X"D3",X"54",X"45",X"50",X"AB",X"AD",X"AA",X"AF",X"DE",X"C1",X"4E",X"44",X"CF",
		X"52",X"BE",X"BD",X"BC",X"D3",X"47",X"4E",X"C9",X"4E",X"54",X"C1",X"42",X"53",X"D5",X"53",X"52",
		X"C6",X"52",X"45",X"CC",X"50",X"4F",X"53",X"D0",X"4F",X"53",X"D3",X"51",X"52",X"D2",X"4E",X"44",
		X"CC",X"4F",X"47",X"C5",X"58",X"50",X"C3",X"4F",X"53",X"D3",X"49",X"4E",X"D4",X"41",X"4E",X"C1",
		X"54",X"4E",X"D0",X"45",X"45",X"4B",X"CC",X"45",X"4E",X"D3",X"54",X"52",X"24",X"D6",X"41",X"4C",
		X"C1",X"53",X"43",X"C3",X"48",X"52",X"24",X"CC",X"45",X"46",X"54",X"24",X"D2",X"49",X"47",X"48",
		X"54",X"24",X"CD",X"49",X"44",X"24",X"D0",X"4F",X"49",X"4E",X"54",X"80",X"79",X"5C",X"16",X"79",
		X"5C",X"12",X"7C",X"C9",X"13",X"7C",X"2D",X"14",X"7F",X"7E",X"17",X"50",X"A9",X"0A",X"46",X"A8",
		X"0A",X"20",X"45",X"72",X"72",X"6F",X"72",X"07",X"00",X"20",X"69",X"6E",X"20",X"00",X"4F",X"6B",
		X"0D",X"0A",X"00",X"42",X"72",X"65",X"61",X"6B",X"00",X"4E",X"46",X"53",X"4E",X"52",X"47",X"4F",
		X"44",X"46",X"43",X"4F",X"56",X"4F",X"4D",X"55",X"4C",X"42",X"53",X"44",X"44",X"2F",X"30",X"49",
		X"44",X"54",X"4D",X"4F",X"53",X"4C",X"53",X"53",X"54",X"43",X"4E",X"55",X"46",X"4D",X"4F",X"21",
		X"04",X"00",X"39",X"7E",X"23",X"FE",X"81",X"C0",X"4E",X"23",X"46",X"23",X"E5",X"60",X"69",X"7A",
		X"B3",X"EB",X"28",X"02",X"EB",X"E7",X"01",X"0D",X"00",X"E1",X"C8",X"09",X"18",X"E5",X"2A",X"C9",
		X"38",X"22",X"4D",X"38",X"1E",X"02",X"01",X"1E",X"14",X"01",X"1E",X"00",X"01",X"1E",X"12",X"01",
		X"1E",X"22",X"01",X"1E",X"0A",X"01",X"1E",X"24",X"01",X"1E",X"18",X"CD",X"E5",X"0B",X"F7",X"00",
		X"CD",X"DE",X"19",X"21",X"79",X"03",X"F7",X"01",X"57",X"19",X"3E",X"3F",X"DF",X"7E",X"DF",X"D7",
		X"DF",X"21",X"61",X"03",X"CD",X"9D",X"0E",X"2A",X"4D",X"38",X"7C",X"A5",X"3C",X"C4",X"6D",X"16",
		X"3E",X"C1",X"F7",X"02",X"CD",X"BE",X"19",X"AF",X"32",X"08",X"38",X"CD",X"DE",X"19",X"21",X"6E",
		X"03",X"CD",X"9D",X"0E",X"21",X"FF",X"FF",X"22",X"4D",X"38",X"CD",X"85",X"0D",X"38",X"F5",X"D7",
		X"3C",X"3D",X"28",X"F0",X"F5",X"CD",X"9C",X"06",X"D5",X"CD",X"BC",X"04",X"47",X"D1",X"F1",X"F7",
		X"03",X"D2",X"4B",X"06",X"D5",X"C5",X"AF",X"32",X"CC",X"38",X"D7",X"B7",X"F5",X"CD",X"9F",X"04",
		X"38",X"06",X"F1",X"F5",X"CA",X"F3",X"06",X"B7",X"C5",X"30",X"10",X"EB",X"2A",X"D6",X"38",X"1A",
		X"02",X"03",X"13",X"E7",X"20",X"F9",X"60",X"69",X"22",X"D6",X"38",X"D1",X"F1",X"28",X"21",X"2A",
		X"D6",X"38",X"E3",X"C1",X"09",X"E5",X"CD",X"92",X"0B",X"E1",X"22",X"D6",X"38",X"EB",X"74",X"D1",
		X"23",X"23",X"73",X"23",X"72",X"23",X"11",X"60",X"38",X"1A",X"77",X"23",X"13",X"B7",X"20",X"F9",
		X"F7",X"04",X"CD",X"CB",X"0B",X"F7",X"05",X"23",X"EB",X"62",X"6B",X"7E",X"23",X"B6",X"CA",X"14",
		X"04",X"23",X"23",X"23",X"AF",X"BE",X"23",X"20",X"FC",X"EB",X"73",X"23",X"72",X"18",X"EA",X"2A",
		X"4F",X"38",X"44",X"4D",X"7E",X"23",X"B6",X"2B",X"C8",X"23",X"23",X"7E",X"23",X"66",X"6F",X"E7",
		X"60",X"69",X"7E",X"23",X"66",X"6F",X"3F",X"C8",X"3F",X"D0",X"18",X"E6",X"AF",X"32",X"AC",X"38",
		X"0E",X"05",X"11",X"60",X"38",X"7E",X"FE",X"20",X"CA",X"3C",X"05",X"47",X"FE",X"22",X"CA",X"58",
		X"05",X"B7",X"CA",X"5E",X"05",X"3A",X"AC",X"38",X"B7",X"7E",X"C2",X"3C",X"05",X"FE",X"3F",X"3E",
		X"95",X"CA",X"3C",X"05",X"7E",X"FE",X"30",X"38",X"05",X"FE",X"3C",X"DA",X"3C",X"05",X"D5",X"11",
		X"44",X"02",X"C5",X"01",X"36",X"05",X"C5",X"06",X"7F",X"7E",X"FE",X"61",X"38",X"07",X"FE",X"7B",
		X"30",X"03",X"E6",X"5F",X"77",X"4E",X"EB",X"23",X"B6",X"F2",X"07",X"05",X"04",X"7E",X"E6",X"7F",
		X"C8",X"B9",X"20",X"F3",X"EB",X"E5",X"13",X"1A",X"B7",X"FA",X"32",X"05",X"4F",X"78",X"FE",X"88",
		X"20",X"02",X"D7",X"2B",X"23",X"7E",X"FE",X"61",X"38",X"02",X"E6",X"5F",X"B9",X"28",X"E7",X"E1",
		X"18",X"D3",X"48",X"F1",X"EB",X"C9",X"F7",X"0A",X"EB",X"79",X"C1",X"D1",X"23",X"12",X"13",X"0C",
		X"D6",X"3A",X"28",X"04",X"FE",X"49",X"20",X"03",X"32",X"AC",X"38",X"D6",X"54",X"C2",X"C5",X"04",
		X"47",X"7E",X"B7",X"28",X"09",X"B8",X"28",X"E4",X"23",X"12",X"0C",X"13",X"18",X"F3",X"21",X"5F",
		X"38",X"12",X"13",X"12",X"13",X"12",X"C9",X"3E",X"01",X"32",X"47",X"38",X"3E",X"17",X"32",X"08",
		X"38",X"CD",X"9C",X"06",X"C0",X"C1",X"CD",X"9F",X"04",X"C5",X"E1",X"4E",X"23",X"46",X"23",X"78",
		X"B1",X"CA",X"02",X"04",X"CD",X"25",X"1A",X"C5",X"CD",X"EA",X"19",X"5E",X"23",X"56",X"23",X"E5",
		X"EB",X"CD",X"75",X"16",X"3E",X"20",X"E1",X"DF",X"7E",X"23",X"B7",X"28",X"DD",X"F2",X"97",X"05",
		X"F7",X"16",X"D6",X"7F",X"4F",X"11",X"45",X"02",X"1A",X"13",X"B7",X"F2",X"A8",X"05",X"0D",X"20",
		X"F7",X"E6",X"7F",X"DF",X"1A",X"13",X"B7",X"F2",X"B1",X"05",X"18",X"DC",X"3E",X"64",X"32",X"CB",
		X"38",X"CD",X"31",X"07",X"C1",X"E5",X"CD",X"1C",X"07",X"22",X"C7",X"38",X"21",X"02",X"00",X"39",
		X"CD",X"A3",X"03",X"20",X"14",X"09",X"D5",X"2B",X"56",X"2B",X"5E",X"23",X"23",X"E5",X"2A",X"C7",
		X"38",X"E7",X"E1",X"D1",X"20",X"EA",X"D1",X"F9",X"0C",X"D1",X"EB",X"0E",X"08",X"CD",X"A0",X"0B",
		X"E5",X"2A",X"C7",X"38",X"E3",X"E5",X"2A",X"4D",X"38",X"E3",X"CD",X"75",X"09",X"CF",X"A1",X"CD",
		X"72",X"09",X"E5",X"CD",X"2E",X"15",X"E1",X"C5",X"D5",X"01",X"00",X"81",X"51",X"5A",X"7E",X"FE",
		X"A7",X"3E",X"01",X"20",X"0A",X"D7",X"CD",X"72",X"09",X"E5",X"CD",X"2E",X"15",X"EF",X"E1",X"C5",
		X"D5",X"F5",X"33",X"E5",X"2A",X"CE",X"38",X"E3",X"06",X"81",X"C5",X"33",X"22",X"CE",X"38",X"CD",
		X"C2",X"1F",X"7E",X"FE",X"3A",X"28",X"14",X"B7",X"C2",X"C4",X"03",X"23",X"7E",X"23",X"B6",X"CA",
		X"29",X"0C",X"23",X"5E",X"23",X"56",X"EB",X"22",X"4D",X"38",X"EB",X"D7",X"11",X"2C",X"06",X"D5",
		X"C8",X"D6",X"80",X"DA",X"31",X"07",X"FE",X"20",X"F7",X"17",X"D2",X"C4",X"03",X"07",X"4F",X"06",
		X"00",X"EB",X"21",X"D5",X"01",X"09",X"4E",X"23",X"46",X"C5",X"EB",X"23",X"7E",X"FE",X"3A",X"D0",
		X"FE",X"20",X"28",X"F7",X"FE",X"30",X"3F",X"3C",X"3D",X"C9",X"D7",X"CD",X"72",X"09",X"EF",X"FA",
		X"97",X"06",X"3A",X"E7",X"38",X"FE",X"90",X"DA",X"86",X"15",X"01",X"80",X"90",X"11",X"00",X"00",
		X"E5",X"CD",X"5B",X"15",X"E1",X"51",X"C8",X"1E",X"08",X"C3",X"DB",X"03",X"2B",X"11",X"00",X"00",
		X"D7",X"D0",X"E5",X"F5",X"21",X"98",X"19",X"E7",X"38",X"11",X"62",X"6B",X"19",X"29",X"19",X"29",
		X"F1",X"D6",X"30",X"5F",X"16",X"00",X"19",X"EB",X"E1",X"18",X"E5",X"F1",X"E1",X"C9",X"F7",X"18",
		X"CA",X"CB",X"0B",X"CD",X"CF",X"0B",X"01",X"2C",X"06",X"18",X"10",X"0E",X"03",X"CD",X"A0",X"0B",
		X"C1",X"E5",X"E5",X"2A",X"4D",X"38",X"E3",X"3E",X"8C",X"F5",X"33",X"C5",X"CD",X"9C",X"06",X"CD",
		X"1E",X"07",X"23",X"E5",X"2A",X"4D",X"38",X"E7",X"E1",X"DC",X"A2",X"04",X"D4",X"9F",X"04",X"60",
		X"69",X"2B",X"D8",X"1E",X"0E",X"C3",X"DB",X"03",X"C0",X"16",X"FF",X"CD",X"9F",X"03",X"F9",X"FE",
		X"8C",X"1E",X"04",X"C2",X"DB",X"03",X"E1",X"22",X"4D",X"38",X"23",X"7C",X"B5",X"20",X"07",X"3A",
		X"CC",X"38",X"B7",X"C2",X"01",X"04",X"21",X"2C",X"06",X"E3",X"3E",X"E1",X"01",X"3A",X"0E",X"00",
		X"06",X"00",X"79",X"48",X"47",X"7E",X"B7",X"C8",X"B8",X"C8",X"23",X"FE",X"22",X"28",X"F3",X"18",
		X"F4",X"CD",X"D1",X"10",X"CF",X"B0",X"D5",X"3A",X"AB",X"38",X"F5",X"CD",X"85",X"09",X"F1",X"E3",
		X"22",X"CE",X"38",X"1F",X"CD",X"77",X"09",X"CA",X"79",X"07",X"E5",X"2A",X"E4",X"38",X"E5",X"23",
		X"23",X"5E",X"23",X"56",X"2A",X"4F",X"38",X"E7",X"30",X"0E",X"2A",X"DA",X"38",X"E7",X"D1",X"30",
		X"0F",X"21",X"BD",X"38",X"E7",X"30",X"09",X"3E",X"D1",X"CD",X"E4",X"0F",X"EB",X"CD",X"39",X"0E",
		X"CD",X"E4",X"0F",X"E1",X"CD",X"3D",X"15",X"E1",X"C9",X"E5",X"CD",X"3A",X"15",X"D1",X"E1",X"C9",
		X"F7",X"19",X"CD",X"54",X"0B",X"7E",X"47",X"FE",X"8C",X"28",X"03",X"CF",X"88",X"2B",X"4B",X"0D",
		X"78",X"CA",X"51",X"06",X"CD",X"9D",X"06",X"FE",X"2C",X"C0",X"18",X"F3",X"CD",X"85",X"09",X"7E",
		X"FE",X"88",X"28",X"03",X"CF",X"A5",X"2B",X"CD",X"75",X"09",X"EF",X"CA",X"1E",X"07",X"D7",X"DA",
		X"DC",X"06",X"C3",X"50",X"06",X"3E",X"01",X"32",X"47",X"38",X"2B",X"D7",X"F7",X"06",X"CC",X"EA",
		X"19",X"CA",X"66",X"08",X"FE",X"A0",X"CA",X"3A",X"08",X"FE",X"A3",X"CA",X"3A",X"08",X"E5",X"FE",
		X"2C",X"28",X"44",X"FE",X"3B",X"CA",X"61",X"08",X"C1",X"CD",X"85",X"09",X"E5",X"3A",X"AB",X"38",
		X"B7",X"C2",X"11",X"08",X"CD",X"80",X"16",X"CD",X"5F",X"0E",X"36",X"20",X"2A",X"E4",X"38",X"3A",
		X"47",X"38",X"B7",X"28",X"08",X"3A",X"46",X"38",X"86",X"FE",X"84",X"18",X"0D",X"3A",X"48",X"38",
		X"47",X"3C",X"28",X"09",X"3A",X"00",X"38",X"86",X"3D",X"B8",X"D4",X"EA",X"19",X"CD",X"A0",X"0E",
		X"AF",X"C4",X"A0",X"0E",X"E1",X"18",X"A3",X"3A",X"47",X"38",X"B7",X"28",X"08",X"3A",X"46",X"38",
		X"FE",X"70",X"C3",X"2D",X"08",X"3A",X"49",X"38",X"47",X"3A",X"00",X"38",X"B8",X"D4",X"EA",X"19",
		X"D2",X"61",X"08",X"D6",X"0E",X"30",X"FC",X"2F",X"18",X"20",X"F5",X"CD",X"53",X"0B",X"CF",X"29",
		X"2B",X"F1",X"D6",X"A3",X"E5",X"28",X"0F",X"3A",X"47",X"38",X"B7",X"CA",X"53",X"08",X"3A",X"46",
		X"38",X"18",X"03",X"3A",X"00",X"38",X"2F",X"83",X"30",X"07",X"3C",X"47",X"3E",X"20",X"DF",X"10",
		X"FD",X"E1",X"D7",X"C3",X"C1",X"07",X"F7",X"07",X"AF",X"32",X"47",X"38",X"C9",X"3F",X"52",X"65",
		X"64",X"6F",X"20",X"66",X"72",X"6F",X"6D",X"20",X"73",X"74",X"61",X"72",X"74",X"0D",X"0A",X"00",
		X"F7",X"08",X"3A",X"CD",X"38",X"B7",X"C2",X"BE",X"03",X"C1",X"21",X"6D",X"08",X"CD",X"9D",X"0E",
		X"C3",X"01",X"0C",X"F7",X"1A",X"CD",X"45",X"0B",X"7E",X"FE",X"22",X"3E",X"00",X"C2",X"AA",X"08",
		X"CD",X"60",X"0E",X"CF",X"3B",X"E5",X"CD",X"A0",X"0E",X"3E",X"E5",X"CD",X"5B",X"0D",X"C1",X"DA",
		X"26",X"0C",X"23",X"7E",X"B7",X"2B",X"C5",X"CA",X"1B",X"07",X"36",X"2C",X"18",X"05",X"E5",X"2A",
		X"DC",X"38",X"F6",X"AF",X"32",X"CD",X"38",X"E3",X"01",X"CF",X"2C",X"CD",X"D1",X"10",X"E3",X"D5",
		X"7E",X"FE",X"2C",X"28",X"1B",X"3A",X"CD",X"38",X"B7",X"C2",X"53",X"09",X"3E",X"3F",X"DF",X"CD",
		X"5B",X"0D",X"D1",X"C1",X"DA",X"26",X"0C",X"23",X"7E",X"2B",X"B7",X"C5",X"CA",X"1B",X"07",X"D5",
		X"F7",X"1C",X"3A",X"AB",X"38",X"B7",X"28",X"1F",X"D7",X"57",X"47",X"FE",X"22",X"28",X"0C",X"3A",
		X"CD",X"38",X"B7",X"57",X"28",X"02",X"16",X"3A",X"06",X"2C",X"2B",X"CD",X"63",X"0E",X"EB",X"21",
		X"20",X"09",X"E3",X"D5",X"C3",X"4A",X"07",X"D7",X"CD",X"E5",X"15",X"E3",X"CD",X"3A",X"15",X"E1",
		X"2B",X"D7",X"28",X"05",X"FE",X"2C",X"C2",X"80",X"08",X"E3",X"2B",X"D7",X"C2",X"C9",X"08",X"D1",
		X"3A",X"CD",X"38",X"B7",X"EB",X"C2",X"1A",X"0C",X"D5",X"B6",X"21",X"42",X"09",X"C4",X"9D",X"0E",
		X"E1",X"C9",X"3F",X"45",X"78",X"74",X"72",X"61",X"20",X"69",X"67",X"6E",X"6F",X"72",X"65",X"64",
		X"0D",X"0A",X"00",X"CD",X"1C",X"07",X"B7",X"20",X"11",X"23",X"7E",X"23",X"B6",X"1E",X"06",X"CA",
		X"DB",X"03",X"23",X"5E",X"23",X"56",X"ED",X"53",X"C9",X"38",X"D7",X"FE",X"83",X"20",X"E4",X"C3",
		X"F0",X"08",X"CD",X"85",X"09",X"F6",X"37",X"3A",X"AB",X"38",X"8F",X"B7",X"E8",X"C3",X"D9",X"03",
		X"CF",X"B0",X"01",X"CF",X"28",X"2B",X"16",X"00",X"D5",X"0E",X"01",X"CD",X"A0",X"0B",X"CD",X"FD",
		X"09",X"22",X"D0",X"38",X"2A",X"D0",X"38",X"C1",X"78",X"FE",X"78",X"D4",X"75",X"09",X"7E",X"22",
		X"C3",X"38",X"FE",X"A8",X"D8",X"FE",X"B2",X"D0",X"FE",X"AF",X"D2",X"E2",X"09",X"D6",X"A8",X"5F",
		X"20",X"08",X"3A",X"AB",X"38",X"3D",X"7B",X"CA",X"7C",X"0F",X"07",X"83",X"5F",X"21",X"4C",X"03",
		X"16",X"00",X"19",X"78",X"56",X"BA",X"D0",X"23",X"CD",X"75",X"09",X"C5",X"01",X"94",X"09",X"C5",
		X"43",X"4A",X"CD",X"13",X"15",X"58",X"51",X"4E",X"23",X"46",X"23",X"C5",X"2A",X"C3",X"38",X"C3",
		X"88",X"09",X"16",X"00",X"D6",X"AF",X"DA",X"D0",X"0A",X"FE",X"03",X"D2",X"D0",X"0A",X"FE",X"01",
		X"17",X"AA",X"BA",X"57",X"DA",X"C4",X"03",X"22",X"C3",X"38",X"D7",X"18",X"E7",X"F7",X"09",X"AF",
		X"32",X"AB",X"38",X"D7",X"CA",X"D6",X"03",X"DA",X"E5",X"15",X"CD",X"C6",X"0C",X"D2",X"4E",X"0A",
		X"FE",X"A8",X"28",X"E9",X"FE",X"2E",X"CA",X"E5",X"15",X"FE",X"A9",X"CA",X"3D",X"0A",X"FE",X"22",
		X"CA",X"60",X"0E",X"FE",X"A6",X"CA",X"05",X"0B",X"FE",X"A4",X"CA",X"FB",X"19",X"FE",X"A2",X"CA",
		X"40",X"0B",X"D6",X"B2",X"D2",X"5F",X"0A",X"CD",X"83",X"09",X"CF",X"29",X"C9",X"16",X"7D",X"CD",
		X"88",X"09",X"2A",X"D0",X"38",X"E5",X"CD",X"0B",X"15",X"CD",X"75",X"09",X"E1",X"C9",X"CD",X"D1",
		X"10",X"E5",X"EB",X"22",X"E4",X"38",X"3A",X"AB",X"38",X"B7",X"CC",X"20",X"15",X"E1",X"C9",X"F7",
		X"1B",X"FE",X"18",X"CA",X"68",X"1A",X"06",X"00",X"07",X"4F",X"C5",X"D7",X"79",X"FE",X"29",X"38",
		X"16",X"CD",X"83",X"09",X"CF",X"2C",X"CD",X"76",X"09",X"EB",X"2A",X"E4",X"38",X"E3",X"E5",X"EB",
		X"CD",X"54",X"0B",X"EB",X"E3",X"18",X"08",X"CD",X"37",X"0A",X"E3",X"11",X"49",X"0A",X"D5",X"01",
		X"15",X"02",X"09",X"4E",X"23",X"66",X"69",X"E9",X"15",X"FE",X"A9",X"C8",X"FE",X"2D",X"C8",X"14",
		X"FE",X"2B",X"C8",X"FE",X"A8",X"C8",X"2B",X"C9",X"F6",X"AF",X"F5",X"CD",X"75",X"09",X"CD",X"82",
		X"06",X"F1",X"EB",X"C1",X"E3",X"EB",X"CD",X"23",X"15",X"F5",X"CD",X"82",X"06",X"F1",X"C1",X"79",
		X"21",X"21",X"0B",X"C2",X"CB",X"0A",X"A3",X"4F",X"78",X"A2",X"E9",X"B3",X"4F",X"78",X"B2",X"E9",
		X"21",X"E2",X"0A",X"3A",X"AB",X"38",X"1F",X"7A",X"17",X"5F",X"16",X"64",X"78",X"BA",X"D0",X"C3",
		X"CB",X"09",X"E4",X"0A",X"79",X"B7",X"1F",X"C1",X"D1",X"F5",X"CD",X"77",X"09",X"21",X"FB",X"0A",
		X"E5",X"CA",X"5B",X"15",X"AF",X"32",X"AB",X"38",X"C3",X"FC",X"0D",X"3C",X"8F",X"C1",X"A0",X"C6",
		X"FF",X"9F",X"C3",X"F6",X"14",X"16",X"5A",X"CD",X"88",X"09",X"CD",X"75",X"09",X"CD",X"82",X"06",
		X"7B",X"2F",X"4F",X"7A",X"2F",X"CD",X"21",X"0B",X"C1",X"C3",X"94",X"09",X"7D",X"93",X"4F",X"7C",
		X"9A",X"41",X"50",X"1E",X"00",X"21",X"AB",X"38",X"73",X"06",X"90",X"C3",X"FB",X"14",X"3A",X"46",
		X"38",X"18",X"03",X"3A",X"00",X"38",X"47",X"AF",X"C3",X"22",X"0B",X"F7",X"0F",X"C3",X"C4",X"03",
		X"F7",X"10",X"C3",X"C4",X"03",X"E5",X"2A",X"4D",X"38",X"23",X"7C",X"B5",X"E1",X"C0",X"1E",X"16",
		X"C3",X"DB",X"03",X"D7",X"CD",X"72",X"09",X"CD",X"7E",X"06",X"7A",X"B7",X"C2",X"97",X"06",X"2B",
		X"D7",X"7B",X"C9",X"CD",X"82",X"06",X"CD",X"88",X"0B",X"1A",X"C3",X"36",X"0B",X"CD",X"72",X"09",
		X"CD",X"82",X"06",X"CD",X"88",X"0B",X"D5",X"CF",X"2C",X"CD",X"54",X"0B",X"D1",X"12",X"C9",X"CD",
		X"85",X"09",X"E5",X"CD",X"82",X"06",X"E1",X"C9",X"E5",X"21",X"FF",X"2F",X"E7",X"E1",X"D2",X"97",
		X"06",X"C9",X"CD",X"A9",X"0B",X"C5",X"E3",X"C1",X"E7",X"7E",X"02",X"C8",X"0B",X"2B",X"18",X"F8",
		X"E5",X"2A",X"DA",X"38",X"06",X"00",X"09",X"09",X"3E",X"E5",X"3E",X"D0",X"95",X"6F",X"3E",X"FF",
		X"9C",X"67",X"38",X"03",X"39",X"E1",X"D8",X"11",X"0C",X"00",X"C3",X"DB",X"03",X"C0",X"F7",X"0C",
		X"2A",X"4F",X"38",X"AF",X"77",X"23",X"77",X"23",X"22",X"D6",X"38",X"2A",X"4F",X"38",X"2B",X"22",
		X"CE",X"38",X"2A",X"AD",X"38",X"22",X"C1",X"38",X"AF",X"CD",X"05",X"0C",X"2A",X"D6",X"38",X"22",
		X"D8",X"38",X"22",X"DA",X"38",X"C1",X"2A",X"4B",X"38",X"F9",X"CD",X"D8",X"1F",X"22",X"AF",X"38",
		X"CD",X"BE",X"19",X"AF",X"6F",X"67",X"22",X"D4",X"38",X"32",X"CB",X"38",X"22",X"DE",X"38",X"E5",
		X"C5",X"2A",X"CE",X"38",X"C9",X"EB",X"2A",X"4F",X"38",X"28",X"0E",X"EB",X"CD",X"9C",X"06",X"E5",
		X"CD",X"9F",X"04",X"60",X"69",X"D1",X"D2",X"F3",X"06",X"2B",X"22",X"DC",X"38",X"EB",X"C9",X"C0",
		X"F6",X"C0",X"22",X"CE",X"38",X"21",X"F6",X"FF",X"C1",X"2A",X"4D",X"38",X"F5",X"7D",X"A4",X"3C",
		X"28",X"09",X"22",X"D2",X"38",X"2A",X"CE",X"38",X"22",X"D4",X"38",X"CD",X"BE",X"19",X"CD",X"DE",
		X"19",X"F1",X"21",X"73",X"03",X"C2",X"F4",X"03",X"C3",X"02",X"04",X"2A",X"D4",X"38",X"7C",X"B5",
		X"11",X"20",X"00",X"CA",X"DB",X"03",X"ED",X"5B",X"D2",X"38",X"ED",X"53",X"4D",X"38",X"C9",X"C3",
		X"97",X"06",X"3E",X"AF",X"B7",X"F5",X"D7",X"3E",X"01",X"32",X"CB",X"38",X"CD",X"D1",X"10",X"C2",
		X"97",X"06",X"32",X"CB",X"38",X"CD",X"75",X"09",X"F1",X"E5",X"F5",X"C5",X"06",X"23",X"28",X"12",
		X"CD",X"7F",X"1B",X"CD",X"BC",X"1B",X"78",X"CD",X"87",X"1B",X"CD",X"87",X"1B",X"CD",X"87",X"1B",
		X"18",X"11",X"CD",X"2E",X"1B",X"CD",X"CE",X"1B",X"0E",X"06",X"CD",X"4D",X"1B",X"B8",X"20",X"F8",
		X"0D",X"20",X"F7",X"E1",X"EB",X"19",X"EB",X"4E",X"06",X"00",X"09",X"09",X"23",X"E7",X"28",X"0D",
		X"F1",X"F5",X"7E",X"C4",X"8A",X"1B",X"CC",X"4D",X"1B",X"77",X"23",X"18",X"F0",X"F1",X"C2",X"1C",
		X"1C",X"E1",X"C3",X"7E",X"1B",X"7E",X"FE",X"41",X"D8",X"FE",X"5B",X"3F",X"C9",X"F7",X"0B",X"CA",
		X"CF",X"0B",X"CD",X"7B",X"06",X"2B",X"D7",X"E5",X"2A",X"AD",X"38",X"28",X"0E",X"E1",X"CF",X"2C",
		X"D5",X"CD",X"7B",X"06",X"2B",X"D7",X"C2",X"C4",X"03",X"E3",X"EB",X"7D",X"93",X"5F",X"7C",X"9A",
		X"57",X"DA",X"B7",X"0B",X"E5",X"2A",X"D6",X"38",X"01",X"28",X"00",X"09",X"E7",X"D2",X"B7",X"0B",
		X"EB",X"22",X"4B",X"38",X"E1",X"22",X"AD",X"38",X"E1",X"C3",X"CF",X"0B",X"7D",X"93",X"5F",X"7C",
		X"9A",X"57",X"C9",X"11",X"00",X"00",X"C4",X"D1",X"10",X"22",X"CE",X"38",X"CD",X"9F",X"03",X"C2",
		X"CA",X"03",X"F9",X"D5",X"7E",X"F5",X"23",X"D5",X"CD",X"20",X"15",X"E3",X"E5",X"CD",X"53",X"12",
		X"E1",X"CD",X"3A",X"15",X"E1",X"CD",X"31",X"15",X"E5",X"CD",X"5B",X"15",X"E1",X"C1",X"90",X"CD",
		X"31",X"15",X"28",X"09",X"EB",X"22",X"4D",X"38",X"69",X"60",X"C3",X"28",X"06",X"F9",X"2A",X"CE",
		X"38",X"7E",X"FE",X"2C",X"C2",X"2C",X"06",X"D7",X"CD",X"16",X"0D",X"3E",X"3F",X"DF",X"3E",X"20",
		X"DF",X"C3",X"85",X"0D",X"3A",X"4A",X"38",X"B7",X"3E",X"5C",X"32",X"4A",X"38",X"20",X"05",X"05",
		X"28",X"13",X"DF",X"04",X"05",X"2B",X"28",X"09",X"7E",X"DF",X"18",X"12",X"05",X"2B",X"DF",X"20",
		X"0D",X"DF",X"CD",X"EA",X"19",X"21",X"60",X"38",X"06",X"01",X"AF",X"32",X"4A",X"38",X"CD",X"DA",
		X"19",X"4F",X"FE",X"7F",X"28",X"CE",X"3A",X"4A",X"38",X"B7",X"28",X"07",X"3E",X"5C",X"DF",X"AF",
		X"32",X"4A",X"38",X"79",X"FE",X"07",X"28",X"41",X"FE",X"03",X"CC",X"EA",X"19",X"37",X"C8",X"FE",
		X"0D",X"CA",X"E5",X"19",X"FE",X"15",X"CA",X"82",X"0D",X"00",X"00",X"00",X"00",X"00",X"FE",X"08",
		X"CA",X"7C",X"0D",X"FE",X"18",X"20",X"05",X"3E",X"23",X"C3",X"81",X"0D",X"FE",X"12",X"20",X"14",
		X"C5",X"D5",X"E5",X"36",X"00",X"CD",X"EA",X"19",X"21",X"60",X"38",X"CD",X"9D",X"0E",X"E1",X"D1",
		X"C1",X"C3",X"8E",X"0D",X"FE",X"20",X"DA",X"8E",X"0D",X"78",X"FE",X"49",X"3E",X"07",X"D2",X"F8",
		X"0D",X"79",X"71",X"32",X"CC",X"38",X"23",X"04",X"DF",X"C3",X"8E",X"0D",X"D5",X"CD",X"C9",X"0F",
		X"7E",X"23",X"23",X"4E",X"23",X"46",X"D1",X"C5",X"F5",X"CD",X"CD",X"0F",X"CD",X"31",X"15",X"F1",
		X"57",X"E1",X"7B",X"B2",X"C8",X"7A",X"D6",X"01",X"D8",X"AF",X"BB",X"3C",X"D0",X"15",X"1D",X"0A",
		X"03",X"BE",X"23",X"28",X"ED",X"3F",X"C3",X"F1",X"14",X"CD",X"75",X"09",X"CD",X"80",X"16",X"CD",
		X"5F",X"0E",X"CD",X"C9",X"0F",X"01",X"1D",X"10",X"C5",X"7E",X"23",X"23",X"E5",X"CD",X"B3",X"0E",
		X"E1",X"4E",X"23",X"46",X"CD",X"53",X"0E",X"E5",X"6F",X"CD",X"BD",X"0F",X"D1",X"C9",X"3E",X"01",
		X"CD",X"B3",X"0E",X"21",X"BD",X"38",X"E5",X"77",X"23",X"23",X"73",X"23",X"72",X"E1",X"C9",X"2B",
		X"06",X"22",X"50",X"E5",X"0E",X"FF",X"23",X"7E",X"0C",X"B7",X"28",X"06",X"BA",X"28",X"03",X"B8",
		X"20",X"F4",X"FE",X"22",X"CC",X"6B",X"06",X"E3",X"23",X"EB",X"79",X"CD",X"53",X"0E",X"11",X"BD",
		X"38",X"2A",X"AF",X"38",X"22",X"E4",X"38",X"3E",X"01",X"32",X"AB",X"38",X"CD",X"3D",X"15",X"E7",
		X"22",X"AF",X"38",X"E1",X"7E",X"C0",X"11",X"1E",X"00",X"C3",X"DB",X"03",X"23",X"CD",X"5F",X"0E",
		X"CD",X"C9",X"0F",X"CD",X"31",X"15",X"1C",X"1D",X"C8",X"0A",X"DF",X"FE",X"0D",X"CC",X"F0",X"19",
		X"03",X"18",X"F4",X"B7",X"0E",X"F1",X"F5",X"2A",X"4B",X"38",X"EB",X"2A",X"C1",X"38",X"2F",X"4F",
		X"06",X"FF",X"09",X"23",X"E7",X"38",X"07",X"22",X"C1",X"38",X"23",X"EB",X"F1",X"C9",X"F1",X"11",
		X"1A",X"00",X"CA",X"DB",X"03",X"BF",X"F5",X"01",X"B5",X"0E",X"C5",X"2A",X"AD",X"38",X"22",X"C1",
		X"38",X"21",X"00",X"00",X"E5",X"2A",X"DA",X"38",X"E5",X"21",X"B1",X"38",X"ED",X"5B",X"AF",X"38",
		X"E7",X"01",X"EC",X"0E",X"C2",X"32",X"0F",X"2A",X"D6",X"38",X"ED",X"5B",X"D8",X"38",X"E7",X"28",
		X"0A",X"23",X"7E",X"23",X"B7",X"CD",X"35",X"0F",X"18",X"F0",X"C1",X"ED",X"5B",X"DA",X"38",X"E7",
		X"CA",X"57",X"0F",X"CD",X"31",X"15",X"7A",X"E5",X"09",X"B7",X"F2",X"0A",X"0F",X"22",X"C5",X"38",
		X"E1",X"4E",X"06",X"00",X"09",X"09",X"23",X"EB",X"2A",X"C5",X"38",X"EB",X"E7",X"28",X"DC",X"01",
		X"27",X"0F",X"C5",X"F6",X"80",X"7E",X"23",X"23",X"5E",X"23",X"56",X"23",X"F0",X"B7",X"C8",X"44",
		X"4D",X"2A",X"C1",X"38",X"E7",X"60",X"69",X"D8",X"E1",X"E3",X"E7",X"E3",X"E5",X"60",X"69",X"D0",
		X"C1",X"F1",X"F1",X"E5",X"D5",X"C5",X"C9",X"D1",X"E1",X"7C",X"B5",X"C8",X"2B",X"46",X"2B",X"4E",
		X"E5",X"2B",X"2B",X"6E",X"26",X"00",X"09",X"50",X"59",X"2B",X"44",X"4D",X"2A",X"C1",X"38",X"CD",
		X"95",X"0B",X"E1",X"71",X"23",X"70",X"60",X"69",X"2B",X"C3",X"DE",X"0E",X"C5",X"E5",X"2A",X"E4",
		X"38",X"E3",X"CD",X"FD",X"09",X"E3",X"CD",X"76",X"09",X"7E",X"E5",X"2A",X"E4",X"38",X"E5",X"86",
		X"11",X"1C",X"00",X"DA",X"DB",X"03",X"CD",X"50",X"0E",X"D1",X"CD",X"CD",X"0F",X"E3",X"CD",X"CC",
		X"0F",X"E5",X"2A",X"BF",X"38",X"EB",X"CD",X"B4",X"0F",X"CD",X"B4",X"0F",X"21",X"91",X"09",X"E3",
		X"E5",X"C3",X"7E",X"0E",X"E1",X"E3",X"7E",X"23",X"23",X"4E",X"23",X"46",X"6F",X"2C",X"2D",X"C8",
		X"0A",X"12",X"03",X"13",X"18",X"F8",X"CD",X"76",X"09",X"2A",X"E4",X"38",X"EB",X"CD",X"E4",X"0F",
		X"EB",X"C0",X"D5",X"50",X"59",X"1B",X"4E",X"2A",X"C1",X"38",X"E7",X"20",X"05",X"47",X"09",X"22",
		X"C1",X"38",X"E1",X"C9",X"2A",X"AF",X"38",X"2B",X"46",X"2B",X"4E",X"2B",X"2B",X"E7",X"C0",X"22",
		X"AF",X"38",X"C9",X"01",X"36",X"0B",X"C5",X"CD",X"C6",X"0F",X"AF",X"57",X"32",X"AB",X"38",X"7E",
		X"B7",X"C9",X"01",X"36",X"0B",X"C5",X"CD",X"F7",X"0F",X"CA",X"97",X"06",X"23",X"23",X"5E",X"23",
		X"56",X"1A",X"C9",X"CD",X"4E",X"0E",X"CD",X"57",X"0B",X"2A",X"BF",X"38",X"73",X"C1",X"C3",X"7E",
		X"0E",X"CD",X"A0",X"10",X"AF",X"E3",X"4F",X"E5",X"7E",X"B8",X"38",X"02",X"78",X"11",X"0E",X"00",
		X"C5",X"CD",X"B3",X"0E",X"C1",X"E1",X"E5",X"23",X"23",X"46",X"23",X"66",X"68",X"06",X"00",X"09",
		X"44",X"4D",X"CD",X"53",X"0E",X"6F",X"CD",X"BD",X"0F",X"D1",X"CD",X"CD",X"0F",X"C3",X"7E",X"0E",
		X"CD",X"A0",X"10",X"D1",X"D5",X"1A",X"90",X"18",X"CC",X"EB",X"7E",X"CD",X"A3",X"10",X"04",X"05",
		X"CA",X"97",X"06",X"C5",X"1E",X"FF",X"FE",X"29",X"28",X"05",X"CF",X"2C",X"CD",X"54",X"0B",X"CF",
		X"29",X"F1",X"E3",X"01",X"27",X"10",X"C5",X"3D",X"BE",X"06",X"00",X"D0",X"4F",X"7E",X"91",X"BB",
		X"47",X"D8",X"43",X"C9",X"CD",X"F7",X"0F",X"CA",X"C3",X"12",X"5F",X"23",X"23",X"7E",X"23",X"66",
		X"6F",X"E5",X"19",X"46",X"72",X"E3",X"C5",X"2B",X"D7",X"CD",X"E5",X"15",X"C1",X"E1",X"70",X"C9",
		X"EB",X"CF",X"29",X"C1",X"D1",X"C5",X"43",X"C9",X"2A",X"DA",X"38",X"EB",X"21",X"00",X"00",X"39",
		X"3A",X"AB",X"38",X"B7",X"CA",X"1C",X"0B",X"CD",X"C9",X"0F",X"CD",X"DB",X"0E",X"ED",X"5B",X"4B",
		X"38",X"2A",X"C1",X"38",X"C3",X"1C",X"0B",X"2B",X"D7",X"C8",X"CF",X"2C",X"01",X"C7",X"10",X"C5",
		X"F6",X"AF",X"32",X"AA",X"38",X"4E",X"CD",X"C5",X"0C",X"DA",X"C4",X"03",X"AF",X"47",X"32",X"AB",
		X"38",X"D7",X"38",X"05",X"CD",X"C6",X"0C",X"38",X"09",X"47",X"D7",X"38",X"FD",X"CD",X"C6",X"0C",
		X"30",X"F8",X"D6",X"24",X"20",X"08",X"3C",X"32",X"AB",X"38",X"0F",X"80",X"47",X"D7",X"3A",X"CB",
		X"38",X"3D",X"CA",X"A0",X"11",X"F2",X"0E",X"11",X"7E",X"D6",X"28",X"CA",X"7A",X"11",X"AF",X"32",
		X"CB",X"38",X"E5",X"50",X"59",X"2A",X"DE",X"38",X"E7",X"11",X"E0",X"38",X"CA",X"1A",X"14",X"2A",
		X"D8",X"38",X"EB",X"2A",X"D6",X"38",X"E7",X"CA",X"3D",X"11",X"79",X"96",X"23",X"C2",X"32",X"11",
		X"78",X"96",X"23",X"CA",X"6C",X"11",X"23",X"23",X"23",X"23",X"C3",X"26",X"11",X"E1",X"E3",X"D5",
		X"11",X"51",X"0A",X"E7",X"D1",X"CA",X"6F",X"11",X"E3",X"E5",X"C5",X"01",X"06",X"00",X"2A",X"DA",
		X"38",X"E5",X"09",X"C1",X"E5",X"CD",X"92",X"0B",X"E1",X"22",X"DA",X"38",X"60",X"69",X"22",X"D8",
		X"38",X"2B",X"36",X"00",X"E7",X"20",X"FA",X"D1",X"73",X"23",X"72",X"23",X"EB",X"E1",X"C9",X"32",
		X"E7",X"38",X"21",X"6D",X"03",X"22",X"E4",X"38",X"E1",X"C9",X"E5",X"2A",X"AA",X"38",X"E3",X"57",
		X"D5",X"C5",X"CD",X"7A",X"06",X"C1",X"F1",X"EB",X"E3",X"E5",X"EB",X"3C",X"57",X"7E",X"FE",X"2C",
		X"CA",X"80",X"11",X"CF",X"29",X"22",X"D0",X"38",X"E1",X"22",X"AA",X"38",X"1E",X"00",X"D5",X"11",
		X"E5",X"F5",X"2A",X"D8",X"38",X"3E",X"19",X"ED",X"5B",X"DA",X"38",X"E7",X"28",X"25",X"7E",X"23",
		X"B9",X"20",X"02",X"7E",X"B8",X"23",X"5E",X"23",X"56",X"23",X"20",X"EA",X"3A",X"AA",X"38",X"B7",
		X"C2",X"CD",X"03",X"F1",X"44",X"4D",X"CA",X"1A",X"14",X"96",X"CA",X"2B",X"12",X"11",X"10",X"00",
		X"C3",X"DB",X"03",X"11",X"04",X"00",X"F1",X"CA",X"97",X"06",X"71",X"23",X"70",X"23",X"4F",X"CD",
		X"A0",X"0B",X"23",X"23",X"22",X"C3",X"38",X"71",X"23",X"3A",X"AA",X"38",X"17",X"79",X"01",X"0B",
		X"00",X"30",X"02",X"C1",X"03",X"71",X"F5",X"23",X"70",X"23",X"E5",X"CD",X"CA",X"15",X"EB",X"E1",
		X"F1",X"3D",X"20",X"EA",X"F5",X"42",X"4B",X"EB",X"19",X"DA",X"B7",X"0B",X"CD",X"A9",X"0B",X"22",
		X"DA",X"38",X"2B",X"36",X"00",X"E7",X"20",X"FA",X"03",X"57",X"2A",X"C3",X"38",X"5E",X"EB",X"29",
		X"09",X"EB",X"2B",X"2B",X"73",X"23",X"72",X"23",X"F1",X"38",X"21",X"47",X"4F",X"7E",X"23",X"16",
		X"E1",X"5E",X"23",X"56",X"23",X"E3",X"F5",X"E7",X"D2",X"CD",X"11",X"E5",X"CD",X"CA",X"15",X"D1",
		X"19",X"F1",X"3D",X"44",X"4D",X"20",X"E9",X"29",X"29",X"C1",X"09",X"EB",X"2A",X"D0",X"38",X"C9",
		X"21",X"57",X"17",X"CD",X"31",X"15",X"18",X"09",X"CD",X"31",X"15",X"21",X"C1",X"D1",X"CD",X"0B",
		X"15",X"78",X"B7",X"C8",X"3A",X"E7",X"38",X"B7",X"CA",X"23",X"15",X"90",X"30",X"0C",X"2F",X"3C",
		X"EB",X"CD",X"13",X"15",X"EB",X"CD",X"23",X"15",X"C1",X"D1",X"FE",X"19",X"D0",X"F5",X"CD",X"46",
		X"15",X"67",X"F1",X"CD",X"30",X"13",X"7C",X"B7",X"21",X"E4",X"38",X"F2",X"9F",X"12",X"CD",X"10",
		X"13",X"30",X"5E",X"23",X"34",X"CA",X"D3",X"03",X"2E",X"01",X"CD",X"52",X"13",X"18",X"52",X"AF",
		X"90",X"47",X"7E",X"9B",X"5F",X"23",X"7E",X"9A",X"57",X"23",X"7E",X"99",X"4F",X"DC",X"1C",X"13",
		X"68",X"63",X"AF",X"47",X"79",X"B7",X"20",X"27",X"4A",X"54",X"65",X"6F",X"78",X"D6",X"08",X"FE",
		X"E0",X"20",X"F0",X"AF",X"32",X"E7",X"38",X"C9",X"7C",X"B5",X"B2",X"20",X"0A",X"79",X"05",X"17",
		X"30",X"FC",X"04",X"1F",X"4F",X"18",X"0B",X"05",X"29",X"7A",X"17",X"57",X"79",X"8F",X"4F",X"F2",
		X"C8",X"12",X"78",X"5C",X"45",X"B7",X"28",X"09",X"21",X"E7",X"38",X"86",X"77",X"30",X"D4",X"28",
		X"D2",X"78",X"21",X"E7",X"38",X"B7",X"FC",X"03",X"13",X"46",X"23",X"7E",X"E6",X"80",X"A9",X"4F",
		X"C3",X"23",X"15",X"1C",X"C0",X"14",X"C0",X"0C",X"C0",X"0E",X"80",X"34",X"C0",X"C3",X"D3",X"03",
		X"7E",X"83",X"5F",X"23",X"7E",X"8A",X"57",X"23",X"7E",X"89",X"4F",X"C9",X"21",X"E8",X"38",X"7E",
		X"2F",X"77",X"AF",X"6F",X"90",X"47",X"7D",X"9B",X"5F",X"7D",X"9A",X"57",X"7D",X"99",X"4F",X"C9",
		X"06",X"00",X"D6",X"08",X"38",X"07",X"43",X"5A",X"51",X"0E",X"00",X"18",X"F5",X"C6",X"09",X"6F",
		X"7A",X"B3",X"B0",X"20",X"09",X"79",X"2D",X"C8",X"1F",X"4F",X"30",X"FA",X"18",X"06",X"AF",X"2D",
		X"C8",X"79",X"1F",X"4F",X"7A",X"1F",X"57",X"7B",X"1F",X"5F",X"78",X"1F",X"47",X"18",X"EF",X"00",
		X"00",X"00",X"81",X"04",X"9A",X"F7",X"19",X"83",X"24",X"63",X"43",X"83",X"75",X"CD",X"8D",X"84",
		X"A9",X"7F",X"83",X"82",X"04",X"00",X"00",X"00",X"81",X"E2",X"B0",X"4D",X"83",X"0A",X"72",X"11",
		X"83",X"F4",X"04",X"35",X"7F",X"EF",X"B7",X"EA",X"97",X"06",X"CD",X"95",X"13",X"01",X"31",X"80",
		X"11",X"18",X"72",X"18",X"36",X"CD",X"2E",X"15",X"3E",X"80",X"32",X"E7",X"38",X"A8",X"F5",X"CD",
		X"13",X"15",X"21",X"63",X"13",X"CD",X"46",X"18",X"C1",X"E1",X"CD",X"13",X"15",X"EB",X"CD",X"23",
		X"15",X"21",X"74",X"13",X"CD",X"46",X"18",X"C1",X"D1",X"CD",X"2F",X"14",X"F1",X"CD",X"13",X"15",
		X"CD",X"F6",X"14",X"C1",X"D1",X"C3",X"61",X"12",X"21",X"C1",X"D1",X"EF",X"C8",X"2E",X"00",X"CD",
		X"AC",X"14",X"79",X"32",X"F6",X"38",X"EB",X"22",X"F7",X"38",X"01",X"00",X"00",X"50",X"58",X"21",
		X"B0",X"12",X"E5",X"21",X"EB",X"13",X"E5",X"E5",X"21",X"E4",X"38",X"7E",X"23",X"B7",X"28",X"2C",
		X"E5",X"2E",X"08",X"1F",X"67",X"79",X"30",X"0B",X"E5",X"2A",X"F7",X"38",X"19",X"EB",X"E1",X"3A",
		X"F6",X"38",X"89",X"1F",X"4F",X"7A",X"1F",X"57",X"7B",X"1F",X"5F",X"78",X"1F",X"47",X"E6",X"10",
		X"28",X"04",X"78",X"F6",X"20",X"47",X"2D",X"7C",X"20",X"D9",X"E1",X"C9",X"43",X"5A",X"51",X"4F",
		X"C9",X"CD",X"13",X"15",X"01",X"20",X"84",X"11",X"00",X"00",X"CD",X"23",X"15",X"C1",X"D1",X"EF",
		X"CA",X"C7",X"03",X"2E",X"FF",X"CD",X"AC",X"14",X"34",X"CA",X"D3",X"03",X"34",X"CA",X"D3",X"03",
		X"2B",X"7E",X"32",X"19",X"38",X"2B",X"7E",X"32",X"15",X"38",X"2B",X"7E",X"32",X"11",X"38",X"41",
		X"EB",X"AF",X"4F",X"57",X"5F",X"32",X"1C",X"38",X"E5",X"C5",X"7D",X"CD",X"10",X"38",X"DE",X"00",
		X"3F",X"30",X"07",X"32",X"1C",X"38",X"F1",X"F1",X"37",X"D2",X"C1",X"E1",X"79",X"3C",X"3D",X"1F",
		X"F2",X"87",X"14",X"17",X"3A",X"1C",X"38",X"1F",X"E6",X"C0",X"F5",X"78",X"B4",X"B5",X"28",X"02",
		X"3E",X"20",X"E1",X"B4",X"C3",X"F2",X"12",X"17",X"7B",X"17",X"5F",X"7A",X"17",X"57",X"79",X"17",
		X"4F",X"29",X"78",X"17",X"47",X"3A",X"1C",X"38",X"17",X"32",X"1C",X"38",X"79",X"B2",X"B3",X"20",
		X"B7",X"E5",X"21",X"E7",X"38",X"35",X"E1",X"20",X"AF",X"C3",X"C3",X"12",X"78",X"B7",X"28",X"1D",
		X"7D",X"21",X"E7",X"38",X"AE",X"80",X"47",X"1F",X"A8",X"78",X"F2",X"CC",X"14",X"C6",X"80",X"77",
		X"CA",X"1A",X"14",X"CD",X"46",X"15",X"77",X"2B",X"C9",X"EF",X"2F",X"E1",X"B7",X"E1",X"F2",X"C3",
		X"12",X"C3",X"D3",X"03",X"CD",X"2E",X"15",X"78",X"B7",X"C8",X"C6",X"02",X"DA",X"D3",X"03",X"47",
		X"CD",X"61",X"12",X"21",X"E7",X"38",X"34",X"C0",X"C3",X"D3",X"03",X"3A",X"E6",X"38",X"FE",X"2F",
		X"17",X"9F",X"C0",X"3C",X"C9",X"EF",X"06",X"88",X"11",X"00",X"00",X"21",X"E7",X"38",X"4F",X"70",
		X"06",X"00",X"23",X"36",X"80",X"17",X"C3",X"AD",X"12",X"EF",X"F0",X"21",X"E6",X"38",X"7E",X"EE",
		X"80",X"77",X"C9",X"EB",X"2A",X"E4",X"38",X"E3",X"E5",X"2A",X"E6",X"38",X"E3",X"E5",X"EB",X"C9",
		X"CD",X"31",X"15",X"EB",X"22",X"E4",X"38",X"60",X"69",X"22",X"E6",X"38",X"EB",X"C9",X"21",X"E4",
		X"38",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"C9",X"11",X"E4",X"38",X"06",X"04",X"1A",
		X"77",X"13",X"23",X"10",X"FA",X"C9",X"21",X"E6",X"38",X"7E",X"07",X"37",X"1F",X"77",X"3F",X"1F",
		X"23",X"23",X"77",X"79",X"07",X"37",X"1F",X"4F",X"1F",X"AE",X"C9",X"78",X"B7",X"CA",X"28",X"00",
		X"21",X"EF",X"14",X"E5",X"EF",X"79",X"C8",X"21",X"E6",X"38",X"AE",X"79",X"F8",X"CD",X"73",X"15",
		X"1F",X"A9",X"C9",X"23",X"78",X"BE",X"C0",X"2B",X"79",X"BE",X"C0",X"2B",X"7A",X"BE",X"C0",X"2B",
		X"7B",X"96",X"C0",X"E1",X"E1",X"C9",X"47",X"4F",X"57",X"5F",X"B7",X"C8",X"E5",X"CD",X"2E",X"15",
		X"CD",X"46",X"15",X"AE",X"67",X"FC",X"AA",X"15",X"3E",X"98",X"90",X"CD",X"30",X"13",X"7C",X"17",
		X"DC",X"03",X"13",X"06",X"00",X"DC",X"1C",X"13",X"E1",X"C9",X"1B",X"7A",X"A3",X"3C",X"C0",X"0B",
		X"C9",X"21",X"E7",X"38",X"7E",X"FE",X"98",X"3A",X"E4",X"38",X"D0",X"7E",X"CD",X"86",X"15",X"36",
		X"98",X"7B",X"F5",X"79",X"17",X"CD",X"AD",X"12",X"F1",X"C9",X"21",X"00",X"00",X"78",X"B1",X"C8",
		X"3E",X"10",X"29",X"DA",X"CD",X"11",X"EB",X"29",X"EB",X"D2",X"E0",X"15",X"09",X"DA",X"CD",X"11",
		X"3D",X"C2",X"D2",X"15",X"C9",X"FE",X"2D",X"F5",X"28",X"05",X"FE",X"2B",X"28",X"01",X"2B",X"CD",
		X"C3",X"12",X"47",X"57",X"5F",X"2F",X"4F",X"D7",X"DA",X"3F",X"16",X"FE",X"2E",X"CA",X"1A",X"16",
		X"FE",X"65",X"CA",X"0A",X"16",X"FE",X"45",X"C2",X"1E",X"16",X"D7",X"CD",X"98",X"0A",X"D7",X"DA",
		X"61",X"16",X"14",X"C2",X"1E",X"16",X"AF",X"93",X"5F",X"0C",X"0C",X"CA",X"F7",X"15",X"E5",X"7B",
		X"90",X"F4",X"37",X"16",X"F2",X"2D",X"16",X"F5",X"CD",X"21",X"14",X"F1",X"3C",X"C2",X"21",X"16",
		X"D1",X"F1",X"CC",X"0B",X"15",X"EB",X"C9",X"C8",X"F5",X"CD",X"D4",X"14",X"F1",X"3D",X"C9",X"D5",
		X"57",X"78",X"89",X"47",X"C5",X"E5",X"D5",X"CD",X"D4",X"14",X"F1",X"D6",X"30",X"CD",X"56",X"16",
		X"E1",X"C1",X"D1",X"C3",X"F7",X"15",X"CD",X"13",X"15",X"CD",X"F6",X"14",X"C1",X"D1",X"C3",X"61",
		X"12",X"7B",X"07",X"07",X"83",X"07",X"86",X"D6",X"30",X"5F",X"C3",X"0E",X"16",X"E5",X"21",X"69",
		X"03",X"CD",X"9D",X"0E",X"E1",X"11",X"9C",X"0E",X"D5",X"EB",X"AF",X"06",X"98",X"CD",X"FB",X"14",
		X"21",X"E9",X"38",X"E5",X"EF",X"36",X"20",X"F2",X"8C",X"16",X"36",X"2D",X"23",X"36",X"30",X"CA",
		X"42",X"17",X"E5",X"FC",X"0B",X"15",X"AF",X"F5",X"CD",X"48",X"17",X"01",X"43",X"91",X"11",X"F8",
		X"4F",X"CD",X"5B",X"15",X"B7",X"E2",X"B9",X"16",X"F1",X"CD",X"38",X"16",X"F5",X"C3",X"9B",X"16",
		X"CD",X"21",X"14",X"F1",X"3C",X"F5",X"CD",X"48",X"17",X"CD",X"50",X"12",X"3C",X"CD",X"86",X"15",
		X"CD",X"23",X"15",X"01",X"06",X"03",X"F1",X"81",X"3C",X"FA",X"D5",X"16",X"FE",X"08",X"D2",X"D5",
		X"16",X"3C",X"47",X"3E",X"02",X"3D",X"3D",X"E1",X"F5",X"11",X"5E",X"17",X"05",X"C2",X"E6",X"16",
		X"36",X"2E",X"23",X"36",X"30",X"23",X"05",X"36",X"2E",X"CC",X"38",X"15",X"C5",X"E5",X"D5",X"CD",
		X"2E",X"15",X"E1",X"06",X"2F",X"04",X"7B",X"96",X"5F",X"23",X"7A",X"9E",X"57",X"23",X"79",X"9E",
		X"4F",X"2B",X"2B",X"D2",X"F5",X"16",X"CD",X"10",X"13",X"23",X"CD",X"23",X"15",X"EB",X"E1",X"70",
		X"23",X"C1",X"0D",X"C2",X"E6",X"16",X"05",X"CA",X"26",X"17",X"2B",X"7E",X"FE",X"30",X"CA",X"1A",
		X"17",X"FE",X"2E",X"C4",X"38",X"15",X"F1",X"CA",X"45",X"17",X"36",X"45",X"23",X"36",X"2B",X"F2",
		X"36",X"17",X"36",X"2D",X"2F",X"3C",X"06",X"2F",X"04",X"D6",X"0A",X"D2",X"38",X"17",X"C6",X"3A",
		X"23",X"70",X"23",X"77",X"23",X"71",X"E1",X"C9",X"01",X"74",X"94",X"11",X"F7",X"23",X"CD",X"5B",
		X"15",X"B7",X"E1",X"E2",X"B0",X"16",X"E9",X"00",X"00",X"00",X"80",X"40",X"42",X"0F",X"A0",X"86",
		X"01",X"10",X"27",X"00",X"E8",X"03",X"00",X"64",X"00",X"00",X"0A",X"00",X"00",X"01",X"00",X"00",
		X"21",X"0B",X"15",X"E3",X"E9",X"CD",X"13",X"15",X"21",X"57",X"17",X"CD",X"20",X"15",X"C1",X"D1",
		X"EF",X"78",X"CA",X"CD",X"17",X"F2",X"8C",X"17",X"B7",X"CA",X"C7",X"03",X"B7",X"CA",X"C4",X"12",
		X"D5",X"C5",X"79",X"F6",X"7F",X"CD",X"2E",X"15",X"F2",X"B5",X"17",X"F5",X"3A",X"E7",X"38",X"FE",
		X"99",X"38",X"03",X"F1",X"18",X"0F",X"F1",X"D5",X"C5",X"CD",X"B1",X"15",X"C1",X"D1",X"F5",X"CD",
		X"5B",X"15",X"E1",X"7C",X"1F",X"E1",X"22",X"E6",X"38",X"E1",X"22",X"E4",X"38",X"DC",X"70",X"17",
		X"CC",X"0B",X"15",X"D5",X"C5",X"CD",X"85",X"13",X"C1",X"D1",X"CD",X"CB",X"13",X"01",X"38",X"81",
		X"11",X"3B",X"AA",X"CD",X"CB",X"13",X"3A",X"E7",X"38",X"FE",X"88",X"30",X"22",X"FE",X"68",X"38",
		X"30",X"CD",X"13",X"15",X"CD",X"B1",X"15",X"C6",X"81",X"C1",X"D1",X"28",X"15",X"F5",X"CD",X"5E",
		X"12",X"21",X"1A",X"18",X"CD",X"46",X"18",X"C1",X"11",X"00",X"00",X"4A",X"C3",X"CB",X"13",X"CD",
		X"13",X"15",X"3A",X"E6",X"38",X"B7",X"F2",X"0E",X"18",X"F1",X"F1",X"C3",X"C3",X"12",X"C3",X"D3",
		X"03",X"01",X"00",X"81",X"11",X"00",X"00",X"C3",X"23",X"15",X"07",X"7C",X"88",X"59",X"74",X"E0",
		X"97",X"26",X"77",X"C4",X"1D",X"1E",X"7A",X"5E",X"50",X"63",X"7C",X"1A",X"FE",X"75",X"7E",X"18",
		X"72",X"31",X"80",X"00",X"00",X"00",X"81",X"CD",X"13",X"15",X"11",X"C9",X"13",X"D5",X"E5",X"CD",
		X"2E",X"15",X"CD",X"CB",X"13",X"E1",X"CD",X"13",X"15",X"7E",X"23",X"CD",X"20",X"15",X"06",X"F1",
		X"C1",X"D1",X"3D",X"C8",X"D5",X"C5",X"F5",X"E5",X"CD",X"CB",X"13",X"E1",X"CD",X"31",X"15",X"E5",
		X"CD",X"61",X"12",X"E1",X"18",X"E9",X"EF",X"21",X"20",X"38",X"FA",X"C4",X"18",X"21",X"41",X"38",
		X"CD",X"20",X"15",X"21",X"20",X"38",X"C8",X"86",X"E6",X"07",X"06",X"00",X"77",X"23",X"87",X"87",
		X"4F",X"09",X"CD",X"31",X"15",X"CD",X"CB",X"13",X"3A",X"1F",X"38",X"3C",X"E6",X"03",X"06",X"00",
		X"FE",X"01",X"88",X"32",X"1F",X"38",X"21",X"C7",X"18",X"87",X"87",X"4F",X"09",X"CD",X"53",X"12",
		X"CD",X"2E",X"15",X"7B",X"59",X"EE",X"4F",X"4F",X"36",X"80",X"2B",X"46",X"36",X"80",X"21",X"1E",
		X"38",X"34",X"7E",X"D6",X"AB",X"20",X"04",X"77",X"0C",X"15",X"1C",X"CD",X"B0",X"12",X"21",X"41",
		X"38",X"C3",X"3A",X"15",X"77",X"2B",X"77",X"2B",X"77",X"18",X"D5",X"68",X"B1",X"46",X"68",X"99",
		X"E9",X"92",X"69",X"10",X"D1",X"75",X"68",X"21",X"53",X"19",X"CD",X"53",X"12",X"3A",X"E7",X"38",
		X"FE",X"77",X"D8",X"3A",X"E6",X"38",X"B7",X"F2",X"F3",X"18",X"E6",X"7F",X"32",X"E6",X"38",X"11",
		X"0B",X"15",X"D5",X"01",X"22",X"7E",X"11",X"83",X"F9",X"CD",X"CB",X"13",X"CD",X"13",X"15",X"CD",
		X"B1",X"15",X"C1",X"D1",X"CD",X"5E",X"12",X"01",X"00",X"7F",X"11",X"00",X"00",X"CD",X"5B",X"15",
		X"FA",X"35",X"19",X"01",X"80",X"7F",X"11",X"00",X"00",X"CD",X"61",X"12",X"01",X"80",X"80",X"11",
		X"00",X"00",X"CD",X"61",X"12",X"EF",X"F4",X"0B",X"15",X"01",X"00",X"7F",X"11",X"00",X"00",X"CD",
		X"61",X"12",X"CD",X"0B",X"15",X"3A",X"E6",X"38",X"B7",X"F5",X"F2",X"42",X"19",X"EE",X"80",X"32",
		X"E6",X"38",X"21",X"5B",X"19",X"CD",X"37",X"18",X"F1",X"F0",X"3A",X"E6",X"38",X"EE",X"80",X"32",
		X"E6",X"38",X"C9",X"DB",X"0F",X"49",X"81",X"00",X"00",X"00",X"7F",X"05",X"FB",X"D7",X"1E",X"86",
		X"65",X"26",X"99",X"87",X"58",X"34",X"23",X"87",X"E1",X"5D",X"A5",X"86",X"DB",X"0F",X"49",X"83",
		X"CD",X"13",X"15",X"CD",X"DD",X"18",X"C1",X"E1",X"CD",X"13",X"15",X"EB",X"CD",X"23",X"15",X"CD",
		X"D7",X"18",X"C3",X"2D",X"14",X"F7",X"0E",X"C3",X"C4",X"03",X"F7",X"0D",X"F5",X"3A",X"47",X"38",
		X"B7",X"CA",X"D6",X"19",X"F1",X"F5",X"FE",X"09",X"20",X"0C",X"3E",X"20",X"DF",X"3A",X"46",X"38",
		X"E6",X"07",X"20",X"F6",X"F1",X"C9",X"F1",X"F5",X"D6",X"0D",X"28",X"0B",X"38",X"0C",X"3A",X"46",
		X"38",X"3C",X"FE",X"84",X"CC",X"C7",X"19",X"32",X"46",X"38",X"F1",X"C3",X"E8",X"1A",X"AF",X"32",
		X"47",X"38",X"3A",X"46",X"38",X"B7",X"C8",X"3E",X"0D",X"CD",X"BB",X"19",X"3E",X"0A",X"CD",X"BB",
		X"19",X"AF",X"32",X"46",X"38",X"C9",X"F1",X"C3",X"72",X"1D",X"CD",X"2F",X"1A",X"C9",X"3A",X"00",
		X"38",X"B7",X"C8",X"18",X"05",X"36",X"00",X"21",X"5F",X"38",X"3E",X"0D",X"DF",X"3E",X"0A",X"DF",
		X"3A",X"47",X"38",X"B7",X"28",X"04",X"AF",X"32",X"46",X"38",X"C9",X"D7",X"E5",X"CD",X"18",X"1A",
		X"28",X"09",X"F5",X"CD",X"4E",X"0E",X"F1",X"5F",X"CD",X"19",X"10",X"21",X"6D",X"03",X"22",X"E4",
		X"38",X"3E",X"01",X"32",X"AB",X"38",X"E1",X"C9",X"E5",X"21",X"0A",X"38",X"7E",X"36",X"00",X"B7",
		X"CC",X"39",X"1A",X"E1",X"C9",X"CD",X"39",X"1A",X"C8",X"32",X"0A",X"38",X"FE",X"13",X"C0",X"AF",
		X"32",X"0A",X"38",X"CD",X"39",X"1A",X"28",X"FB",X"C9",X"CD",X"7E",X"1E",X"FE",X"03",X"20",X"0A",
		X"3A",X"5E",X"38",X"B7",X"CC",X"BE",X"0B",X"C3",X"CE",X"1F",X"B7",X"C9",X"AF",X"18",X"02",X"3E",
		X"01",X"08",X"CD",X"7F",X"1A",X"CD",X"8E",X"1A",X"28",X"02",X"36",X"A0",X"08",X"B7",X"1A",X"20",
		X"03",X"2F",X"A6",X"06",X"B6",X"77",X"E1",X"C9",X"D7",X"CD",X"7F",X"1A",X"CD",X"8E",X"1A",X"20",
		X"06",X"1A",X"A6",X"16",X"01",X"20",X"02",X"16",X"00",X"AF",X"CD",X"23",X"0B",X"E1",X"C9",X"CF",
		X"28",X"CD",X"D0",X"1A",X"D5",X"CF",X"2C",X"CD",X"D0",X"1A",X"CF",X"29",X"C1",X"C9",X"E3",X"E5",
		X"C5",X"D5",X"21",X"47",X"00",X"E7",X"DA",X"97",X"06",X"21",X"4F",X"00",X"C5",X"D1",X"E7",X"38",
		X"F5",X"D1",X"C1",X"21",X"28",X"30",X"7B",X"11",X"28",X"00",X"FE",X"03",X"38",X"06",X"19",X"3D",
		X"3D",X"3D",X"18",X"F6",X"07",X"CB",X"29",X"30",X"01",X"3C",X"09",X"11",X"CA",X"1A",X"B7",X"28",
		X"04",X"13",X"3D",X"18",X"F9",X"7E",X"F6",X"A0",X"AE",X"C9",X"01",X"02",X"04",X"08",X"10",X"40",
		X"CD",X"85",X"09",X"C3",X"82",X"06",X"D5",X"CD",X"7F",X"1A",X"E5",X"CD",X"64",X"1E",X"E1",X"D1",
		X"C9",X"3E",X"0D",X"CD",X"E8",X"1A",X"3E",X"0A",X"F7",X"11",X"F5",X"F5",X"D9",X"DB",X"FE",X"E6",
		X"01",X"28",X"FA",X"CD",X"08",X"1B",X"1E",X"08",X"F1",X"CD",X"0A",X"1B",X"0F",X"1D",X"20",X"F9",
		X"3E",X"01",X"CD",X"0A",X"1B",X"D9",X"F1",X"C9",X"3E",X"00",X"D3",X"FE",X"26",X"B1",X"25",X"20",
		X"FD",X"00",X"00",X"00",X"C9",X"E5",X"D5",X"CD",X"E1",X"1A",X"21",X"28",X"30",X"11",X"E8",X"33",
		X"7E",X"CD",X"E8",X"1A",X"23",X"E7",X"38",X"F8",X"CD",X"E1",X"1A",X"D1",X"E1",X"C9",X"E5",X"D5",
		X"C5",X"21",X"E8",X"1B",X"F5",X"CD",X"9D",X"0E",X"21",X"B5",X"00",X"CD",X"9D",X"0E",X"CD",X"7E",
		X"1E",X"FE",X"0D",X"20",X"F9",X"CD",X"EA",X"19",X"F1",X"C1",X"D1",X"E1",X"C9",X"D9",X"0E",X"FC",
		X"CD",X"62",X"1B",X"38",X"FB",X"26",X"08",X"CD",X"62",X"1B",X"CB",X"15",X"25",X"20",X"F8",X"7D",
		X"D9",X"C9",X"ED",X"78",X"1F",X"38",X"FB",X"ED",X"78",X"1F",X"30",X"FB",X"AF",X"3C",X"ED",X"40",
		X"CB",X"18",X"38",X"F9",X"3C",X"ED",X"40",X"CB",X"18",X"30",X"F9",X"FE",X"49",X"C9",X"C9",X"E5",
		X"D5",X"C5",X"21",X"F7",X"1B",X"18",X"AD",X"CD",X"8A",X"1B",X"F5",X"D9",X"0E",X"FC",X"F5",X"AF",
		X"1E",X"01",X"CD",X"A5",X"1B",X"F1",X"1E",X"08",X"CD",X"A5",X"1B",X"3E",X"FF",X"1E",X"02",X"CD",
		X"A5",X"1B",X"D9",X"F1",X"C9",X"17",X"2E",X"40",X"38",X"02",X"2E",X"80",X"06",X"04",X"ED",X"41",
		X"65",X"25",X"20",X"FD",X"05",X"20",X"F7",X"1D",X"20",X"EB",X"C9",X"C9",X"F5",X"C5",X"06",X"0C",
		X"3E",X"FF",X"CD",X"8A",X"1B",X"10",X"F9",X"AF",X"CD",X"8A",X"1B",X"C1",X"F1",X"C9",X"F5",X"C5",
		X"06",X"06",X"CD",X"4D",X"1B",X"3C",X"20",X"F8",X"10",X"F8",X"CD",X"4D",X"1B",X"B7",X"28",X"05",
		X"3C",X"28",X"F7",X"18",X"EB",X"C1",X"F1",X"C9",X"50",X"72",X"65",X"73",X"73",X"20",X"3C",X"50",
		X"4C",X"41",X"59",X"3E",X"0D",X"0A",X"00",X"50",X"72",X"65",X"73",X"73",X"20",X"3C",X"52",X"45",
		X"43",X"4F",X"52",X"44",X"3E",X"0D",X"0A",X"00",X"F7",X"15",X"FE",X"AA",X"CA",X"62",X"0C",X"CD",
		X"B8",X"1C",X"E5",X"CD",X"25",X"1D",X"2A",X"4F",X"38",X"CD",X"38",X"1D",X"06",X"0F",X"AF",X"CD",
		X"8A",X"1B",X"10",X"FB",X"01",X"40",X"1F",X"CD",X"4B",X"1D",X"E1",X"C9",X"F7",X"14",X"FE",X"AA",
		X"CA",X"63",X"0C",X"D6",X"95",X"28",X"02",X"AF",X"01",X"2F",X"23",X"FE",X"01",X"F5",X"3E",X"FF",
		X"32",X"5E",X"38",X"CD",X"B1",X"1C",X"AF",X"32",X"5D",X"38",X"D5",X"CD",X"2E",X"1B",X"CD",X"D9",
		X"1C",X"21",X"57",X"38",X"CD",X"ED",X"1C",X"D1",X"28",X"12",X"21",X"06",X"1D",X"CD",X"0D",X"1D",
		X"06",X"0A",X"CD",X"4D",X"1B",X"B7",X"20",X"F8",X"10",X"F8",X"18",X"DA",X"21",X"FE",X"1C",X"CD",
		X"0D",X"1D",X"F1",X"32",X"E4",X"38",X"DC",X"BE",X"0B",X"3A",X"E4",X"38",X"FE",X"01",X"32",X"5E",
		X"38",X"2A",X"4F",X"38",X"CD",X"51",X"1D",X"20",X"11",X"22",X"D6",X"38",X"21",X"6E",X"03",X"CD",
		X"9D",X"0E",X"3E",X"FF",X"32",X"5E",X"38",X"C3",X"80",X"04",X"23",X"EB",X"2A",X"D6",X"38",X"E7",
		X"38",X"EA",X"21",X"AB",X"1C",X"CD",X"9D",X"0E",X"C3",X"01",X"04",X"42",X"61",X"64",X"0D",X"0A",
		X"00",X"AF",X"32",X"51",X"38",X"2B",X"D7",X"C8",X"CD",X"85",X"09",X"E5",X"CD",X"06",X"10",X"2B",
		X"2B",X"2B",X"46",X"0E",X"06",X"21",X"51",X"38",X"1A",X"77",X"23",X"13",X"0D",X"28",X"08",X"10",
		X"F7",X"41",X"36",X"00",X"23",X"10",X"FB",X"E1",X"C9",X"CD",X"CE",X"1B",X"AF",X"32",X"5D",X"38",
		X"21",X"57",X"38",X"06",X"06",X"CD",X"4D",X"1B",X"77",X"23",X"10",X"F9",X"C9",X"01",X"51",X"38",
		X"1E",X"06",X"0A",X"B7",X"C8",X"0A",X"BE",X"23",X"03",X"C0",X"1D",X"20",X"F8",X"C9",X"46",X"6F",
		X"75",X"6E",X"64",X"3A",X"20",X"00",X"53",X"6B",X"69",X"70",X"3A",X"20",X"00",X"D5",X"F5",X"CD",
		X"9D",X"0E",X"21",X"57",X"38",X"06",X"06",X"7E",X"23",X"B7",X"28",X"01",X"DF",X"10",X"F8",X"CD",
		X"EA",X"19",X"F1",X"D1",X"C9",X"CD",X"7F",X"1B",X"CD",X"BC",X"1B",X"06",X"06",X"21",X"51",X"38",
		X"7E",X"23",X"CD",X"8A",X"1B",X"10",X"F9",X"C9",X"CD",X"BC",X"1B",X"EB",X"2A",X"D6",X"38",X"1A",
		X"13",X"CD",X"8A",X"1B",X"E7",X"20",X"F8",X"C9",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",
		X"C9",X"CD",X"CE",X"1B",X"3E",X"FF",X"32",X"5D",X"38",X"9F",X"2F",X"57",X"06",X"0A",X"CD",X"4D",
		X"1B",X"5F",X"96",X"A2",X"C0",X"73",X"CD",X"A9",X"0B",X"7E",X"B7",X"23",X"20",X"EE",X"10",X"EE",
		X"AF",X"C9",X"F7",X"13",X"F5",X"FE",X"0A",X"28",X"1A",X"3A",X"00",X"38",X"B7",X"20",X"14",X"3A",
		X"08",X"38",X"B7",X"28",X"0E",X"3D",X"32",X"08",X"38",X"20",X"08",X"3E",X"17",X"32",X"08",X"38",
		X"CD",X"2F",X"1A",X"F1",X"F5",X"D9",X"FE",X"07",X"CA",X"14",X"1E",X"FE",X"0B",X"CA",X"45",X"1E",
		X"5F",X"2A",X"01",X"38",X"3A",X"0D",X"38",X"77",X"7B",X"FE",X"08",X"28",X"30",X"FE",X"0D",X"28",
		X"0D",X"FE",X"0A",X"28",X"13",X"2A",X"01",X"38",X"77",X"CD",X"1F",X"1E",X"18",X"2C",X"ED",X"5B",
		X"00",X"38",X"AF",X"57",X"ED",X"52",X"18",X"1F",X"11",X"C0",X"33",X"E7",X"D2",X"D8",X"1D",X"11",
		X"28",X"00",X"19",X"22",X"01",X"38",X"18",X"12",X"CD",X"FE",X"1D",X"18",X"0D",X"3A",X"00",X"38",
		X"B7",X"28",X"02",X"2B",X"3D",X"36",X"20",X"CD",X"3E",X"1E",X"2A",X"01",X"38",X"7E",X"32",X"0D",
		X"38",X"36",X"7F",X"D9",X"F1",X"C9",X"2A",X"01",X"38",X"3A",X"0D",X"38",X"77",X"C9",X"01",X"98",
		X"03",X"11",X"28",X"30",X"21",X"50",X"30",X"ED",X"B0",X"06",X"28",X"21",X"C1",X"33",X"36",X"20",
		X"23",X"10",X"FB",X"C9",X"01",X"C8",X"00",X"11",X"32",X"00",X"CD",X"64",X"1E",X"18",X"D4",X"2A",
		X"01",X"38",X"3A",X"00",X"38",X"23",X"3C",X"FE",X"26",X"38",X"13",X"23",X"23",X"11",X"E8",X"33",
		X"E7",X"3E",X"00",X"38",X"09",X"21",X"C1",X"33",X"CD",X"3E",X"1E",X"C3",X"FE",X"1D",X"22",X"01",
		X"38",X"32",X"00",X"38",X"C9",X"06",X"20",X"21",X"00",X"30",X"CD",X"59",X"1E",X"06",X"06",X"CD",
		X"59",X"1E",X"21",X"29",X"30",X"AF",X"C3",X"E7",X"1D",X"11",X"FF",X"03",X"70",X"23",X"1B",X"7A",
		X"B3",X"20",X"F9",X"C9",X"78",X"B1",X"C8",X"AF",X"D3",X"FC",X"CD",X"76",X"1E",X"3C",X"D3",X"FC",
		X"CD",X"76",X"1E",X"0B",X"18",X"EE",X"D5",X"E1",X"7C",X"B5",X"C8",X"2B",X"18",X"FA",X"F7",X"12",
		X"D9",X"2A",X"0B",X"38",X"7C",X"B7",X"28",X"1A",X"EB",X"21",X"0F",X"38",X"34",X"7E",X"FE",X"0F",
		X"38",X"3C",X"36",X"05",X"EB",X"23",X"7E",X"22",X"0B",X"38",X"B7",X"F2",X"36",X"1F",X"AF",X"32",
		X"0C",X"38",X"01",X"FF",X"00",X"ED",X"78",X"2F",X"E6",X"3F",X"21",X"0E",X"38",X"28",X"16",X"06",
		X"7F",X"ED",X"78",X"2F",X"E6",X"0F",X"20",X"1F",X"06",X"BF",X"ED",X"78",X"2F",X"E6",X"3F",X"20",
		X"16",X"CB",X"08",X"38",X"F5",X"23",X"3E",X"46",X"BE",X"38",X"03",X"28",X"04",X"34",X"AF",X"D9",
		X"C9",X"34",X"2B",X"36",X"00",X"18",X"F7",X"11",X"00",X"00",X"1C",X"1F",X"30",X"FC",X"7B",X"CB",
		X"18",X"30",X"04",X"C6",X"06",X"18",X"F8",X"5F",X"BE",X"77",X"23",X"20",X"0F",X"3E",X"04",X"BE",
		X"38",X"05",X"28",X"0C",X"34",X"18",X"02",X"36",X"06",X"AF",X"D9",X"C9",X"36",X"00",X"18",X"F9",
		X"34",X"06",X"7F",X"ED",X"78",X"CB",X"6F",X"DD",X"21",X"93",X"1F",X"28",X"0C",X"CB",X"67",X"DD",
		X"21",X"65",X"1F",X"28",X"04",X"DD",X"21",X"37",X"1F",X"DD",X"19",X"DD",X"7E",X"00",X"B7",X"F2",
		X"36",X"1F",X"D6",X"7F",X"4F",X"21",X"44",X"02",X"23",X"7E",X"B7",X"F2",X"28",X"1F",X"0D",X"20",
		X"F7",X"22",X"0B",X"38",X"E6",X"7F",X"D9",X"C9",X"3D",X"08",X"3A",X"0D",X"3B",X"2E",X"2D",X"2F",
		X"30",X"70",X"6C",X"2C",X"39",X"6F",X"6B",X"6D",X"6E",X"6A",X"38",X"69",X"37",X"75",X"68",X"62",
		X"36",X"79",X"67",X"76",X"63",X"66",X"35",X"74",X"34",X"72",X"64",X"78",X"33",X"65",X"73",X"7A",
		X"20",X"61",X"32",X"77",X"31",X"71",X"2B",X"5C",X"2A",X"0D",X"40",X"3E",X"5F",X"5E",X"3F",X"50",
		X"4C",X"3C",X"29",X"4F",X"4B",X"4D",X"4E",X"4A",X"28",X"49",X"27",X"55",X"48",X"42",X"26",X"59",
		X"47",X"56",X"43",X"46",X"25",X"54",X"24",X"52",X"44",X"58",X"23",X"45",X"53",X"5A",X"20",X"41",
		X"22",X"57",X"21",X"51",X"82",X"1C",X"C1",X"0D",X"94",X"C4",X"81",X"1E",X"30",X"10",X"CA",X"C3",
		X"92",X"0F",X"9D",X"0D",X"C8",X"9C",X"8D",X"09",X"8C",X"15",X"08",X"C9",X"90",X"19",X"07",X"C7",
		X"03",X"83",X"88",X"84",X"A5",X"12",X"86",X"18",X"8A",X"85",X"13",X"9A",X"C6",X"9B",X"97",X"8E",
		X"89",X"11",X"E5",X"21",X"04",X"00",X"39",X"22",X"F9",X"38",X"E1",X"C3",X"25",X"1A",X"2A",X"F9",
		X"38",X"F9",X"2A",X"CE",X"38",X"CD",X"20",X"0C",X"2B",X"2B",X"22",X"F9",X"38",X"21",X"B1",X"38",
		X"C9",X"3E",X"FF",X"D3",X"FE",X"C3",X"41",X"00",X"3E",X"AA",X"D3",X"FF",X"32",X"09",X"38",X"C3",
		X"10",X"20",X"21",X"5F",X"01",X"C3",X"9D",X"0E",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5",X"F5");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
