library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity char_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of char_rom is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3C",X"20",X"20",X"78",X"20",X"60",X"AC",X"00",X"44",X"48",X"50",X"2C",X"44",X"08",X"1C",X"00",
		X"44",X"48",X"50",X"2C",X"54",X"1C",X"04",X"00",X"64",X"28",X"50",X"2C",X"54",X"1C",X"04",X"00",
		X"00",X"10",X"00",X"7C",X"00",X"10",X"00",X"00",X"3C",X"42",X"99",X"A1",X"A1",X"99",X"42",X"3C",
		X"00",X"04",X"02",X"FF",X"FF",X"02",X"04",X"00",X"00",X"20",X"40",X"FF",X"FF",X"40",X"20",X"00",
		X"18",X"3C",X"5A",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"5A",X"3C",X"18",
		X"0F",X"07",X"0F",X"1D",X"38",X"70",X"20",X"00",X"00",X"04",X"0E",X"1C",X"B8",X"F0",X"E0",X"F0",
		X"00",X"20",X"70",X"38",X"1D",X"0F",X"07",X"0F",X"F0",X"E0",X"F0",X"B8",X"1C",X"0E",X"04",X"00",
		X"00",X"3C",X"3C",X"00",X"7E",X"FF",X"FF",X"FF",X"FC",X"FC",X"3C",X"30",X"30",X"30",X"30",X"30",
		X"FF",X"3C",X"3C",X"3C",X"3C",X"00",X"00",X"00",X"7F",X"7F",X"78",X"18",X"18",X"18",X"18",X"18",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"00",X"3C",X"3C",X"00",X"7E",X"FF",X"BD",X"DB",
		X"7E",X"3C",X"66",X"66",X"E7",X"C3",X"C3",X"C3",X"00",X"38",X"3C",X"00",X"38",X"78",X"7C",X"7F",
		X"7C",X"3E",X"1B",X"1E",X"1C",X"18",X"38",X"38",X"00",X"38",X"3C",X"00",X"39",X"79",X"DF",X"DC",
		X"7C",X"3F",X"1F",X"3B",X"F3",X"C3",X"80",X"00",X"18",X"3C",X"66",X"24",X"E7",X"BD",X"99",X"DB",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"00",
		X"28",X"28",X"28",X"00",X"00",X"00",X"00",X"00",X"28",X"28",X"7C",X"28",X"7C",X"28",X"28",X"00",
		X"10",X"3C",X"50",X"38",X"14",X"78",X"10",X"00",X"60",X"64",X"08",X"10",X"20",X"4C",X"0C",X"00",
		X"20",X"50",X"50",X"20",X"54",X"48",X"34",X"00",X"08",X"08",X"10",X"00",X"00",X"00",X"00",X"00",
		X"10",X"20",X"40",X"40",X"40",X"20",X"10",X"00",X"10",X"08",X"04",X"04",X"04",X"08",X"10",X"00",
		X"10",X"54",X"38",X"10",X"38",X"54",X"10",X"00",X"00",X"10",X"10",X"7C",X"10",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"7C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"04",X"08",X"10",X"20",X"40",X"00",X"00",
		X"38",X"44",X"4C",X"54",X"64",X"44",X"38",X"00",X"10",X"30",X"10",X"10",X"10",X"10",X"38",X"00",
		X"38",X"44",X"04",X"18",X"20",X"40",X"7C",X"00",X"7C",X"04",X"08",X"18",X"04",X"44",X"38",X"00",
		X"08",X"18",X"28",X"48",X"78",X"08",X"08",X"00",X"7C",X"40",X"78",X"04",X"04",X"44",X"38",X"00",
		X"1C",X"20",X"40",X"78",X"44",X"44",X"38",X"00",X"7C",X"04",X"08",X"10",X"20",X"20",X"20",X"00",
		X"38",X"44",X"44",X"38",X"44",X"44",X"38",X"00",X"38",X"44",X"44",X"3C",X"04",X"08",X"70",X"00",
		X"00",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"10",X"10",X"20",X"00",
		X"08",X"10",X"20",X"40",X"20",X"10",X"08",X"00",X"00",X"00",X"7C",X"00",X"7C",X"00",X"00",X"00",
		X"20",X"10",X"08",X"04",X"08",X"10",X"20",X"00",X"38",X"44",X"08",X"10",X"10",X"00",X"10",X"00",
		X"38",X"44",X"54",X"5C",X"58",X"40",X"38",X"00",X"10",X"28",X"44",X"44",X"7C",X"44",X"44",X"00",
		X"78",X"44",X"44",X"78",X"44",X"44",X"78",X"00",X"38",X"44",X"40",X"40",X"40",X"44",X"38",X"00",
		X"78",X"44",X"44",X"44",X"44",X"44",X"78",X"00",X"7C",X"40",X"40",X"78",X"40",X"40",X"7C",X"00",
		X"7C",X"40",X"40",X"78",X"40",X"40",X"40",X"00",X"3C",X"40",X"40",X"40",X"4C",X"44",X"3C",X"00",
		X"44",X"44",X"44",X"7C",X"44",X"44",X"44",X"00",X"38",X"10",X"10",X"10",X"10",X"10",X"38",X"00",
		X"04",X"04",X"04",X"04",X"04",X"44",X"38",X"00",X"44",X"48",X"50",X"60",X"50",X"48",X"44",X"00",
		X"40",X"40",X"40",X"40",X"40",X"40",X"7C",X"00",X"44",X"6C",X"54",X"54",X"44",X"44",X"44",X"00",
		X"44",X"44",X"64",X"54",X"4C",X"44",X"44",X"00",X"38",X"44",X"44",X"44",X"44",X"44",X"38",X"00",
		X"78",X"44",X"44",X"78",X"40",X"40",X"40",X"00",X"38",X"44",X"44",X"44",X"54",X"48",X"34",X"00",
		X"78",X"44",X"44",X"78",X"50",X"48",X"44",X"00",X"38",X"44",X"40",X"38",X"04",X"44",X"38",X"00",
		X"7C",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"44",X"44",X"44",X"44",X"44",X"44",X"38",X"00",
		X"44",X"44",X"44",X"44",X"44",X"28",X"10",X"00",X"44",X"44",X"44",X"54",X"54",X"6C",X"44",X"00",
		X"44",X"44",X"28",X"10",X"28",X"44",X"44",X"00",X"44",X"44",X"28",X"10",X"10",X"10",X"10",X"00",
		X"7C",X"04",X"08",X"10",X"20",X"40",X"7C",X"00",X"7C",X"60",X"60",X"60",X"60",X"60",X"7C",X"00",
		X"00",X"40",X"20",X"10",X"08",X"04",X"00",X"00",X"7C",X"0C",X"0C",X"0C",X"0C",X"0C",X"7C",X"00",
		X"00",X"00",X"10",X"28",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",
		X"20",X"20",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"4C",X"44",X"4C",X"34",X"00",
		X"40",X"40",X"58",X"64",X"44",X"64",X"58",X"00",X"00",X"00",X"1C",X"20",X"20",X"20",X"1C",X"00",
		X"04",X"04",X"34",X"4C",X"44",X"4C",X"34",X"00",X"00",X"00",X"38",X"44",X"7C",X"40",X"38",X"00",
		X"08",X"10",X"10",X"38",X"10",X"10",X"10",X"00",X"00",X"00",X"34",X"4C",X"44",X"3C",X"04",X"38",
		X"40",X"40",X"78",X"44",X"44",X"44",X"44",X"00",X"10",X"00",X"30",X"10",X"10",X"10",X"38",X"00",
		X"08",X"00",X"08",X"08",X"08",X"08",X"08",X"30",X"40",X"40",X"48",X"50",X"70",X"48",X"44",X"00",
		X"30",X"10",X"10",X"10",X"10",X"10",X"38",X"00",X"00",X"00",X"6C",X"52",X"52",X"52",X"52",X"00",
		X"00",X"00",X"78",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"38",X"44",X"44",X"44",X"38",X"00",
		X"00",X"00",X"58",X"64",X"44",X"64",X"58",X"40",X"00",X"00",X"34",X"4C",X"44",X"4C",X"34",X"06",
		X"00",X"00",X"58",X"60",X"40",X"40",X"40",X"00",X"00",X"00",X"3C",X"40",X"38",X"04",X"78",X"00",
		X"10",X"10",X"7C",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"3C",X"00",
		X"00",X"00",X"44",X"44",X"28",X"28",X"10",X"00",X"00",X"00",X"52",X"52",X"52",X"52",X"2C",X"00",
		X"00",X"00",X"44",X"28",X"10",X"28",X"44",X"00",X"00",X"00",X"24",X"24",X"24",X"3C",X"04",X"38",
		X"00",X"00",X"7C",X"08",X"10",X"20",X"7C",X"00",X"0C",X"10",X"10",X"20",X"10",X"10",X"0C",X"00",
		X"10",X"10",X"10",X"00",X"10",X"10",X"10",X"00",X"60",X"10",X"10",X"08",X"10",X"10",X"60",X"00",
		X"00",X"00",X"04",X"38",X"40",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"1C",X"3C",X"00",X"1C",X"1E",X"3E",X"FE",X"3E",X"7C",X"D8",X"78",X"38",X"18",X"1C",X"1C",
		X"00",X"00",X"00",X"00",X"AA",X"55",X"AA",X"55",X"A0",X"50",X"A0",X"50",X"A0",X"50",X"A0",X"50",
		X"AA",X"55",X"AA",X"55",X"AA",X"55",X"AA",X"55",X"00",X"18",X"3C",X"7E",X"7E",X"3C",X"18",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"18",X"3C",X"7E",X"FF",X"DB",X"18",X"3C",X"3C",X"18",X"DB",X"FF",X"7E",X"3C",X"18",X"18",
		X"00",X"1C",X"3C",X"00",X"9C",X"9E",X"FB",X"3B",X"3E",X"FC",X"F8",X"DC",X"CF",X"C3",X"01",X"00",
		X"C0",X"F0",X"FC",X"FF",X"FF",X"FC",X"F0",X"C0",X"18",X"18",X"3C",X"3C",X"7E",X"7E",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"3C",X"52",X"3C",X"80",X"BC",X"FF",X"3D",X"3D",X"3C",X"4A",X"3C",X"01",X"3D",X"FF",X"BC",X"BC",
		X"AA",X"55",X"AA",X"54",X"00",X"00",X"00",X"00",X"0A",X"05",X"0A",X"05",X"0A",X"05",X"0A",X"05",
		X"3C",X"7E",X"FF",X"FF",X"FF",X"FF",X"7E",X"3C",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"30",X"38",X"9C",X"FF",X"FF",X"9C",X"38",X"30",X"0C",X"1C",X"39",X"FF",X"FF",X"39",X"1C",X"0C",
		X"00",X"66",X"7E",X"42",X"C3",X"FF",X"18",X"00",X"00",X"18",X"FF",X"C3",X"42",X"7E",X"66",X"00",
		X"03",X"0F",X"3F",X"FF",X"FF",X"3F",X"0F",X"03",X"FF",X"FF",X"7E",X"7E",X"3C",X"3C",X"18",X"18",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"0F",X"0F",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0F",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"FF",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"00",X"00",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"00",X"00",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",
		X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",
		X"FF",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"00",X"3C",X"3C",X"3C",X"3C",X"00",X"00",X"18",X"3C",X"7E",X"FF",X"FF",X"7E",X"3C",X"18",
		X"00",X"00",X"00",X"18",X"18",X"00",X"00",X"00",X"0F",X"0F",X"07",X"03",X"00",X"00",X"00",X"00",
		X"18",X"18",X"18",X"FF",X"FF",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F0",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"18",X"18",X"18",X"FF",X"FF",X"00",X"00",X"00",X"18",X"18",X"18",X"1F",X"1F",X"18",X"18",X"18",
		X"00",X"00",X"00",X"F8",X"F8",X"18",X"18",X"18",X"18",X"18",X"18",X"1F",X"1F",X"00",X"00",X"00",
		X"09",X"20",X"04",X"80",X"11",X"40",X"08",X"02",X"52",X"44",X"2D",X"C4",X"11",X"B4",X"23",X"4A",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",X"00",X"10",X"2C",X"3A",X"5C",X"34",X"04",X"00",
		X"66",X"FF",X"FF",X"FF",X"7E",X"3C",X"18",X"18",X"18",X"3C",X"18",X"42",X"E7",X"42",X"18",X"3C",
		X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"00",X"00",X"00",X"00",X"03",X"07",X"1F",X"1F",
		X"81",X"42",X"24",X"18",X"18",X"24",X"42",X"81",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",
		X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01",X"C0",X"E0",X"F0",X"F0",X"F0",X"F0",X"E0",X"C0",
		X"00",X"00",X"00",X"FF",X"FF",X"18",X"18",X"18",X"18",X"18",X"18",X"F8",X"F8",X"18",X"18",X"18",
		X"00",X"00",X"00",X"1F",X"1F",X"18",X"18",X"18",X"18",X"18",X"18",X"F8",X"F8",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"F0",X"F0",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"F0",X"F0",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"FF",X"FF",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"00",X"00",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"F0",X"F0",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"0F",X"0F",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
